library ieee;
use ieee.std_logic_1164.all;
use IEEE.Numeric_Std.all;

entity ROMMemory_x16 is
	port(
	address : in  std_logic_vector(15 downto 0);
	data: out std_logic_vector(15 downto 0));
end ROMMemory_x16;

architecture skeleton of ROMMemory_x16 is

	--type rom_array is array (0 to 65535) of std_logic_vector (15 downto 0);
	type rom_array is array (0 to 65535) of std_logic_vector (15 downto 0);
	
	constant rom : rom_array := (
 
  -- Write your algorithm here
  -- :)
	
  -- Início algoritmo que calcula os 20 primeiros números da sequência de Fibonacci
  --0000000000000000 ,  0000000000000001 ,  0000000000000010 ,  0000000000000011 ,  0000000000000100
	"1101001000000001", "1101001010001001", "1101001111111001", "0000101110101000", "1101010000010001", -- 00000 - 00004
	
  --0000000000000101 ,  0000000000000110 ,  0000000000000111 ,  0000000000001000 ,  0000000000001001
	"0101101110000000", "1010000000001111", "1101001100100000", "0100001110101000", "1010000000001100", -- 00005 - 00009
 
  --0000000000001010 ,  0000000000001011 ,  0000000000001100 ,  0000000000001101 ,  0000000000001110
	"1101001100101000", "0100001110001001", "1010000000001001", "1101011000100000", "0000011000101000", -- 00010 - 00014
	
  --0000000000001111 ,  0000000000010000 ,  0000000000010001 ,  0000000000010010 ,  0000000000010011
	"1101001101100000", "1101001000101000", "1101001010110000", "0000110000001000", "0101110000111000", -- 00015 - 00019
  -- Fim algoritmo que calcula os 20 primeiros números da sequência de Fibonacci
  --0000000000010100 ,  0000000000010101 ,  0000000000010110 ,  0000000000010111 ,  0000000000011000
	"1010011111111001", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00020 - 00024
  
  
  
  -- Início algoritmo que calcula os números primos entre 10 e 100
  --0000000000011001 ,  0000000000011010 ,  0000000000011011 ,  0000000000011100 ,  0000000000011101
	"1101001001010001", "1101011001100001", "1101010011101001", "0000010011100000", "0000010011001000", -- 00025 - 00029 
	
  --0000000000011110 ,  0000000000011111 ,  0000000000100000 ,  0000000000100001 ,  0000000000100010
	"0000010011001000", "1101001010100000", "1101001110101000", "1101010000010001", "0111101111000000", -- 00030 - 00034 
 																										
  --0000000000100011 ,  0000000000100100 ,  0000000000100101 ,  0000000000100110 ,  0000000000100111
	"1101001100010000", "0100010000110000", "1010000000000110", "0111101111000000", "0100000010000000", -- 00035 - 00039
	
  --0000000000101000 ,  0000000000101001 ,  0000000000101010 ,  0000000000101011 ,  0000000000101100
	"1010000000000100", "0000110000001000", "1000111111111010", "1101010110111000", "0000101010001000", -- 00040 - 00044 
  -- Fim algoritmo que calcula os números primos entre 10 e 100
  --0000000000101101 ,  0000000000101110 ,  0000000000101111 ,  0000000000110000 ,  0000000000110001
	"0100001011001000", "1010111111110010", "0000000000000000", "0000000000000000", "0000000000000000", -- 00045 - 00049
  
  
  
  -- Início algoritmo que ordena um vetor de 5 posições usando o Bubble Sort
  --0000000000110010 ,  0000000000110011 ,  0000000000110100 ,  0000000000110101 ,  0000000000110110
	"1000100000010001", "1101011010000001", "0100011010101000", "1010000000100000", "1101011110100000", -- 00050 - 00054

  --0000000000110111 ,  0000000000111000 ,  0000000000111001 ,  0000000000111010 ,  0000000000111011
	"0000011111101000", "1011010111111000", "0000111010001000", "1000111111111010", "1101011010000001", -- 00055 - 00059 
	
  --0000000000111100 ,  0000000000111101 ,  0000000000111110 ,  0000000000111111 ,  0000000001000000
	"0100011010101000", "1010000000101110", "1101011110100000", "0000011111101000", "1011010111111000", -- 00060 - 00064 
	
  --0000000001000001 ,  0000000001000010 ,  0000000001000011 ,  0000000001000100 ,  0000000001000101
	"0000111010001000", "1000111111111010", "1101001000000001", "1101001010101001", "1101011000100000", -- 00065 - 00069

  --0000000001000110 ,  0000000001000111 ,  0000000001001000 ,  0000000001001001 ,  0000000001001010
	"1101011010101001", "1100011011100000", "0000111000001000", "1101011010011001", "1100011011100000", -- 00070 - 00074
	
  --0000000001001011 ,  0000000001001100 ,  0000000001001101 ,  0000000001001110 ,  0000000001001111
	"0000111000001000", "1101011011001001", "1100011011100000", "0000111000001000", "1101011010111001", -- 00075 - 00079 
	
  --0000000001010000 ,  0000000001010001 ,  0000000001010010 ,  0000000001010011 ,  0000000001010100
	"1100011011100000", "0000111000001000", "1101011010001001", "1100011011100000", "1000111111011111", -- 00080 - 00084 
	
  --0000000001010101 ,  0000000001010110 ,  0000000001010111 ,  0000000001011000 ,  0000000001011001
	"1101011000000001", "1101011010101000", "0000111010001001", "1101011100000001", "1101011111101000", -- 00085 - 00089
	
  --0000000001011010 ,  0000000001011011 ,  0000000001011100 ,  0000000001011101 ,  0000000001011110
	"0000011111100001", "1101001100100000", "0000001101110000", "1011010110110000", "0000101100001000", -- 00090 - 00094 
	
  --0000000001011111 ,  0000000001100000 ,  0000000001100001 ,  0000000001100010 ,  0000000001100011
	"1011010100110000", "0101010101011000", "1010100000000100", "1100010110110000", "0000101100001001", -- 00095 - 00099
	
  --0000000001100100    0000000001100101    0000000001100110    0000000001100111    0000000001101000  
	"1100010100110000", "0000111100001000", "0101011101111000", "1010011111110100", "0000111000001000", -- 00100 - 00104
  -- Fim algoritmo que ordena um vetor de 5 posições usando o Bubble Sort
  --0000000001101001    0000000001101010    0000000001101011    0000000001101100    0000000001101101
	"0101011001101000", "1010011111101110", "1000111111010000", "0000000000000000", "0000000000000000", -- 00105 - 00109
	
	
	
  -- Espaço não alocado na memória
  --0000000001101110    0000000001101111    0000000001110000    0000000001110001    0000000001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00110 - 00114

  --0000000001110011    0000000001110100    0000000001110101    0000000001110110    0000000001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00115 - 00119

  --0000000001111000    0000000001111001    0000000001111010    0000000001111011    0000000001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00120 - 00124

  --0000000001111101    0000000001111110    0000000001111111    0000000010000000    0000000010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00125 - 00129

  --0000000010000010    0000000010000011    0000000010000100    0000000010000101    0000000010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00130 - 00134

  --0000000010000111    0000000010001000    0000000010001001    0000000010001010    0000000010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00135 - 00139

  --0000000010001100    0000000010001101    0000000010001110    0000000010001111    0000000010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00140 - 00144

  --0000000010010001    0000000010010010    0000000010010011    0000000010010100    0000000010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00145 - 00149

  --0000000010010110    0000000010010111    0000000010011000    0000000010011001    0000000010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00150 - 00154

  --0000000010011011    0000000010011100    0000000010011101    0000000010011110    0000000010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00155 - 00159

  --0000000010100000    0000000010100001    0000000010100010    0000000010100011    0000000010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00160 - 00164

  --0000000010100101    0000000010100110    0000000010100111    0000000010101000    0000000010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00165 - 00169

  --0000000010101010    0000000010101011    0000000010101100    0000000010101101    0000000010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00170 - 00174

  --0000000010101111    0000000010110000    0000000010110001    0000000010110010    0000000010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00175 - 00179

  --0000000010110100    0000000010110101    0000000010110110    0000000010110111    0000000010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00180 - 00184

  --0000000010111001    0000000010111010    0000000010111011    0000000010111100    0000000010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00185 - 00189

  --0000000010111110    0000000010111111    0000000011000000    0000000011000001    0000000011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00190 - 00194

  --0000000011000011    0000000011000100    0000000011000101    0000000011000110    0000000011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00195 - 00199

  --0000000011001000    0000000011001001    0000000011001010    0000000011001011    0000000011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00200 - 00204

  --0000000011001101    0000000011001110    0000000011001111    0000000011010000    0000000011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00205 - 00209

  --0000000011010010    0000000011010011    0000000011010100    0000000011010101    0000000011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00210 - 00214

  --0000000011010111    0000000011011000    0000000011011001    0000000011011010    0000000011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00215 - 00219

  --0000000011011100    0000000011011101    0000000011011110    0000000011011111    0000000011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00220 - 00224

  --0000000011100001    0000000011100010    0000000011100011    0000000011100100    0000000011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00225 - 00229

  --0000000011100110    0000000011100111    0000000011101000    0000000011101001    0000000011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00230 - 00234

  --0000000011101011    0000000011101100    0000000011101101    0000000011101110    0000000011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00235 - 00239

  --0000000011110000    0000000011110001    0000000011110010    0000000011110011    0000000011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00240 - 00244

  --0000000011110101    0000000011110110    0000000011110111    0000000011111000    0000000011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00245 - 00249

  --0000000011111010    0000000011111011    0000000011111100    0000000011111101    0000000011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00250 - 00254

  --0000000011111111    0000000100000000    0000000100000001    0000000100000010    0000000100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00255 - 00259

  --0000000100000100    0000000100000101    0000000100000110    0000000100000111    0000000100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00260 - 00264

  --0000000100001001    0000000100001010    0000000100001011    0000000100001100    0000000100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00265 - 00269

  --0000000100001110    0000000100001111    0000000100010000    0000000100010001    0000000100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00270 - 00274

  --0000000100010011    0000000100010100    0000000100010101    0000000100010110    0000000100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00275 - 00279

  --0000000100011000    0000000100011001    0000000100011010    0000000100011011    0000000100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00280 - 00284

  --0000000100011101    0000000100011110    0000000100011111    0000000100100000    0000000100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00285 - 00289

  --0000000100100010    0000000100100011    0000000100100100    0000000100100101    0000000100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00290 - 00294

  --0000000100100111    0000000100101000    0000000100101001    0000000100101010    0000000100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00295 - 00299

  --0000000100101100    0000000100101101    0000000100101110    0000000100101111    0000000100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00300 - 00304

  --0000000100110001    0000000100110010    0000000100110011    0000000100110100    0000000100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00305 - 00309

  --0000000100110110    0000000100110111    0000000100111000    0000000100111001    0000000100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00310 - 00314

  --0000000100111011    0000000100111100    0000000100111101    0000000100111110    0000000100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00315 - 00319

  --0000000101000000    0000000101000001    0000000101000010    0000000101000011    0000000101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00320 - 00324

  --0000000101000101    0000000101000110    0000000101000111    0000000101001000    0000000101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00325 - 00329

  --0000000101001010    0000000101001011    0000000101001100    0000000101001101    0000000101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00330 - 00334

  --0000000101001111    0000000101010000    0000000101010001    0000000101010010    0000000101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00335 - 00339

  --0000000101010100    0000000101010101    0000000101010110    0000000101010111    0000000101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00340 - 00344

  --0000000101011001    0000000101011010    0000000101011011    0000000101011100    0000000101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00345 - 00349

  --0000000101011110    0000000101011111    0000000101100000    0000000101100001    0000000101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00350 - 00354

  --0000000101100011    0000000101100100    0000000101100101    0000000101100110    0000000101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00355 - 00359

  --0000000101101000    0000000101101001    0000000101101010    0000000101101011    0000000101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00360 - 00364

  --0000000101101101    0000000101101110    0000000101101111    0000000101110000    0000000101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00365 - 00369

  --0000000101110010    0000000101110011    0000000101110100    0000000101110101    0000000101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00370 - 00374

  --0000000101110111    0000000101111000    0000000101111001    0000000101111010    0000000101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00375 - 00379

  --0000000101111100    0000000101111101    0000000101111110    0000000101111111    0000000110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00380 - 00384

  --0000000110000001    0000000110000010    0000000110000011    0000000110000100    0000000110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00385 - 00389

  --0000000110000110    0000000110000111    0000000110001000    0000000110001001    0000000110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00390 - 00394

  --0000000110001011    0000000110001100    0000000110001101    0000000110001110    0000000110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00395 - 00399

  --0000000110010000    0000000110010001    0000000110010010    0000000110010011    0000000110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00400 - 00404

  --0000000110010101    0000000110010110    0000000110010111    0000000110011000    0000000110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00405 - 00409

  --0000000110011010    0000000110011011    0000000110011100    0000000110011101    0000000110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00410 - 00414

  --0000000110011111    0000000110100000    0000000110100001    0000000110100010    0000000110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00415 - 00419

  --0000000110100100    0000000110100101    0000000110100110    0000000110100111    0000000110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00420 - 00424

  --0000000110101001    0000000110101010    0000000110101011    0000000110101100    0000000110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00425 - 00429

  --0000000110101110    0000000110101111    0000000110110000    0000000110110001    0000000110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00430 - 00434

  --0000000110110011    0000000110110100    0000000110110101    0000000110110110    0000000110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00435 - 00439

  --0000000110111000    0000000110111001    0000000110111010    0000000110111011    0000000110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00440 - 00444

  --0000000110111101    0000000110111110    0000000110111111    0000000111000000    0000000111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00445 - 00449

  --0000000111000010    0000000111000011    0000000111000100    0000000111000101    0000000111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00450 - 00454

  --0000000111000111    0000000111001000    0000000111001001    0000000111001010    0000000111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00455 - 00459

  --0000000111001100    0000000111001101    0000000111001110    0000000111001111    0000000111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00460 - 00464

  --0000000111010001    0000000111010010    0000000111010011    0000000111010100    0000000111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00465 - 00469

  --0000000111010110    0000000111010111    0000000111011000    0000000111011001    0000000111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00470 - 00474

  --0000000111011011    0000000111011100    0000000111011101    0000000111011110    0000000111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00475 - 00479

  --0000000111100000    0000000111100001    0000000111100010    0000000111100011    0000000111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00480 - 00484

  --0000000111100101    0000000111100110    0000000111100111    0000000111101000    0000000111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00485 - 00489

  --0000000111101010    0000000111101011    0000000111101100    0000000111101101    0000000111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00490 - 00494

  --0000000111101111    0000000111110000    0000000111110001    0000000111110010    0000000111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00495 - 00499

  --0000000111110100    0000000111110101    0000000111110110    0000000111110111    0000000111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00500 - 00504

  --0000000111111001    0000000111111010    0000000111111011    0000000111111100    0000000111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00505 - 00509

  --0000000111111110    0000000111111111    0000001000000000    0000001000000001    0000001000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00510 - 00514

  --0000001000000011    0000001000000100    0000001000000101    0000001000000110    0000001000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00515 - 00519

  --0000001000001000    0000001000001001    0000001000001010    0000001000001011    0000001000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00520 - 00524

  --0000001000001101    0000001000001110    0000001000001111    0000001000010000    0000001000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00525 - 00529

  --0000001000010010    0000001000010011    0000001000010100    0000001000010101    0000001000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00530 - 00534

  --0000001000010111    0000001000011000    0000001000011001    0000001000011010    0000001000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00535 - 00539

  --0000001000011100    0000001000011101    0000001000011110    0000001000011111    0000001000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00540 - 00544

  --0000001000100001    0000001000100010    0000001000100011    0000001000100100    0000001000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00545 - 00549

  --0000001000100110    0000001000100111    0000001000101000    0000001000101001    0000001000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00550 - 00554

  --0000001000101011    0000001000101100    0000001000101101    0000001000101110    0000001000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00555 - 00559

  --0000001000110000    0000001000110001    0000001000110010    0000001000110011    0000001000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00560 - 00564

  --0000001000110101    0000001000110110    0000001000110111    0000001000111000    0000001000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00565 - 00569

  --0000001000111010    0000001000111011    0000001000111100    0000001000111101    0000001000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00570 - 00574

  --0000001000111111    0000001001000000    0000001001000001    0000001001000010    0000001001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00575 - 00579

  --0000001001000100    0000001001000101    0000001001000110    0000001001000111    0000001001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00580 - 00584

  --0000001001001001    0000001001001010    0000001001001011    0000001001001100    0000001001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00585 - 00589

  --0000001001001110    0000001001001111    0000001001010000    0000001001010001    0000001001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00590 - 00594

  --0000001001010011    0000001001010100    0000001001010101    0000001001010110    0000001001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00595 - 00599

  --0000001001011000    0000001001011001    0000001001011010    0000001001011011    0000001001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00600 - 00604

  --0000001001011101    0000001001011110    0000001001011111    0000001001100000    0000001001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00605 - 00609

  --0000001001100010    0000001001100011    0000001001100100    0000001001100101    0000001001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00610 - 00614

  --0000001001100111    0000001001101000    0000001001101001    0000001001101010    0000001001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00615 - 00619

  --0000001001101100    0000001001101101    0000001001101110    0000001001101111    0000001001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00620 - 00624

  --0000001001110001    0000001001110010    0000001001110011    0000001001110100    0000001001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00625 - 00629

  --0000001001110110    0000001001110111    0000001001111000    0000001001111001    0000001001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00630 - 00634

  --0000001001111011    0000001001111100    0000001001111101    0000001001111110    0000001001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00635 - 00639

  --0000001010000000    0000001010000001    0000001010000010    0000001010000011    0000001010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00640 - 00644

  --0000001010000101    0000001010000110    0000001010000111    0000001010001000    0000001010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00645 - 00649

  --0000001010001010    0000001010001011    0000001010001100    0000001010001101    0000001010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00650 - 00654

  --0000001010001111    0000001010010000    0000001010010001    0000001010010010    0000001010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00655 - 00659

  --0000001010010100    0000001010010101    0000001010010110    0000001010010111    0000001010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00660 - 00664

  --0000001010011001    0000001010011010    0000001010011011    0000001010011100    0000001010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00665 - 00669

  --0000001010011110    0000001010011111    0000001010100000    0000001010100001    0000001010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00670 - 00674

  --0000001010100011    0000001010100100    0000001010100101    0000001010100110    0000001010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00675 - 00679

  --0000001010101000    0000001010101001    0000001010101010    0000001010101011    0000001010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00680 - 00684

  --0000001010101101    0000001010101110    0000001010101111    0000001010110000    0000001010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00685 - 00689

  --0000001010110010    0000001010110011    0000001010110100    0000001010110101    0000001010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00690 - 00694

  --0000001010110111    0000001010111000    0000001010111001    0000001010111010    0000001010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00695 - 00699

  --0000001010111100    0000001010111101    0000001010111110    0000001010111111    0000001011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00700 - 00704

  --0000001011000001    0000001011000010    0000001011000011    0000001011000100    0000001011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00705 - 00709

  --0000001011000110    0000001011000111    0000001011001000    0000001011001001    0000001011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00710 - 00714

  --0000001011001011    0000001011001100    0000001011001101    0000001011001110    0000001011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00715 - 00719

  --0000001011010000    0000001011010001    0000001011010010    0000001011010011    0000001011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00720 - 00724

  --0000001011010101    0000001011010110    0000001011010111    0000001011011000    0000001011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00725 - 00729

  --0000001011011010    0000001011011011    0000001011011100    0000001011011101    0000001011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00730 - 00734

  --0000001011011111    0000001011100000    0000001011100001    0000001011100010    0000001011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00735 - 00739

  --0000001011100100    0000001011100101    0000001011100110    0000001011100111    0000001011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00740 - 00744

  --0000001011101001    0000001011101010    0000001011101011    0000001011101100    0000001011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00745 - 00749

  --0000001011101110    0000001011101111    0000001011110000    0000001011110001    0000001011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00750 - 00754

  --0000001011110011    0000001011110100    0000001011110101    0000001011110110    0000001011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00755 - 00759

  --0000001011111000    0000001011111001    0000001011111010    0000001011111011    0000001011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00760 - 00764

  --0000001011111101    0000001011111110    0000001011111111    0000001100000000    0000001100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00765 - 00769

  --0000001100000010    0000001100000011    0000001100000100    0000001100000101    0000001100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00770 - 00774

  --0000001100000111    0000001100001000    0000001100001001    0000001100001010    0000001100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00775 - 00779

  --0000001100001100    0000001100001101    0000001100001110    0000001100001111    0000001100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00780 - 00784

  --0000001100010001    0000001100010010    0000001100010011    0000001100010100    0000001100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00785 - 00789

  --0000001100010110    0000001100010111    0000001100011000    0000001100011001    0000001100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00790 - 00794

  --0000001100011011    0000001100011100    0000001100011101    0000001100011110    0000001100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00795 - 00799

  --0000001100100000    0000001100100001    0000001100100010    0000001100100011    0000001100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00800 - 00804

  --0000001100100101    0000001100100110    0000001100100111    0000001100101000    0000001100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00805 - 00809

  --0000001100101010    0000001100101011    0000001100101100    0000001100101101    0000001100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00810 - 00814

  --0000001100101111    0000001100110000    0000001100110001    0000001100110010    0000001100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00815 - 00819

  --0000001100110100    0000001100110101    0000001100110110    0000001100110111    0000001100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00820 - 00824

  --0000001100111001    0000001100111010    0000001100111011    0000001100111100    0000001100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00825 - 00829

  --0000001100111110    0000001100111111    0000001101000000    0000001101000001    0000001101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00830 - 00834

  --0000001101000011    0000001101000100    0000001101000101    0000001101000110    0000001101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00835 - 00839

  --0000001101001000    0000001101001001    0000001101001010    0000001101001011    0000001101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00840 - 00844

  --0000001101001101    0000001101001110    0000001101001111    0000001101010000    0000001101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00845 - 00849

  --0000001101010010    0000001101010011    0000001101010100    0000001101010101    0000001101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00850 - 00854

  --0000001101010111    0000001101011000    0000001101011001    0000001101011010    0000001101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00855 - 00859

  --0000001101011100    0000001101011101    0000001101011110    0000001101011111    0000001101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00860 - 00864

  --0000001101100001    0000001101100010    0000001101100011    0000001101100100    0000001101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00865 - 00869

  --0000001101100110    0000001101100111    0000001101101000    0000001101101001    0000001101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00870 - 00874

  --0000001101101011    0000001101101100    0000001101101101    0000001101101110    0000001101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00875 - 00879

  --0000001101110000    0000001101110001    0000001101110010    0000001101110011    0000001101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00880 - 00884

  --0000001101110101    0000001101110110    0000001101110111    0000001101111000    0000001101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00885 - 00889

  --0000001101111010    0000001101111011    0000001101111100    0000001101111101    0000001101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00890 - 00894

  --0000001101111111    0000001110000000    0000001110000001    0000001110000010    0000001110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00895 - 00899

  --0000001110000100    0000001110000101    0000001110000110    0000001110000111    0000001110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00900 - 00904

  --0000001110001001    0000001110001010    0000001110001011    0000001110001100    0000001110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00905 - 00909

  --0000001110001110    0000001110001111    0000001110010000    0000001110010001    0000001110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00910 - 00914

  --0000001110010011    0000001110010100    0000001110010101    0000001110010110    0000001110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00915 - 00919

  --0000001110011000    0000001110011001    0000001110011010    0000001110011011    0000001110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00920 - 00924

  --0000001110011101    0000001110011110    0000001110011111    0000001110100000    0000001110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00925 - 00929

  --0000001110100010    0000001110100011    0000001110100100    0000001110100101    0000001110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00930 - 00934

  --0000001110100111    0000001110101000    0000001110101001    0000001110101010    0000001110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00935 - 00939

  --0000001110101100    0000001110101101    0000001110101110    0000001110101111    0000001110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00940 - 00944

  --0000001110110001    0000001110110010    0000001110110011    0000001110110100    0000001110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00945 - 00949

  --0000001110110110    0000001110110111    0000001110111000    0000001110111001    0000001110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00950 - 00954

  --0000001110111011    0000001110111100    0000001110111101    0000001110111110    0000001110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00955 - 00959

  --0000001111000000    0000001111000001    0000001111000010    0000001111000011    0000001111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00960 - 00964

  --0000001111000101    0000001111000110    0000001111000111    0000001111001000    0000001111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00965 - 00969

  --0000001111001010    0000001111001011    0000001111001100    0000001111001101    0000001111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00970 - 00974

  --0000001111001111    0000001111010000    0000001111010001    0000001111010010    0000001111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00975 - 00979

  --0000001111010100    0000001111010101    0000001111010110    0000001111010111    0000001111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00980 - 00984

  --0000001111011001    0000001111011010    0000001111011011    0000001111011100    0000001111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00985 - 00989

  --0000001111011110    0000001111011111    0000001111100000    0000001111100001    0000001111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00990 - 00994

  --0000001111100011    0000001111100100    0000001111100101    0000001111100110    0000001111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 00995 - 00999

  --0000001111101000    0000001111101001    0000001111101010    0000001111101011    0000001111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01000 - 01004

  --0000001111101101    0000001111101110    0000001111101111    0000001111110000    0000001111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01005 - 01009

  --0000001111110010    0000001111110011    0000001111110100    0000001111110101    0000001111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01010 - 01014

  --0000001111110111    0000001111111000    0000001111111001    0000001111111010    0000001111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01015 - 01019

  --0000001111111100    0000001111111101    0000001111111110    0000001111111111    0000010000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01020 - 01024

  --0000010000000001    0000010000000010    0000010000000011    0000010000000100    0000010000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01025 - 01029

  --0000010000000110    0000010000000111    0000010000001000    0000010000001001    0000010000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01030 - 01034

  --0000010000001011    0000010000001100    0000010000001101    0000010000001110    0000010000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01035 - 01039

  --0000010000010000    0000010000010001    0000010000010010    0000010000010011    0000010000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01040 - 01044

  --0000010000010101    0000010000010110    0000010000010111    0000010000011000    0000010000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01045 - 01049

  --0000010000011010    0000010000011011    0000010000011100    0000010000011101    0000010000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01050 - 01054

  --0000010000011111    0000010000100000    0000010000100001    0000010000100010    0000010000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01055 - 01059

  --0000010000100100    0000010000100101    0000010000100110    0000010000100111    0000010000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01060 - 01064

  --0000010000101001    0000010000101010    0000010000101011    0000010000101100    0000010000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01065 - 01069

  --0000010000101110    0000010000101111    0000010000110000    0000010000110001    0000010000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01070 - 01074

  --0000010000110011    0000010000110100    0000010000110101    0000010000110110    0000010000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01075 - 01079

  --0000010000111000    0000010000111001    0000010000111010    0000010000111011    0000010000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01080 - 01084

  --0000010000111101    0000010000111110    0000010000111111    0000010001000000    0000010001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01085 - 01089

  --0000010001000010    0000010001000011    0000010001000100    0000010001000101    0000010001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01090 - 01094

  --0000010001000111    0000010001001000    0000010001001001    0000010001001010    0000010001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01095 - 01099

  --0000010001001100    0000010001001101    0000010001001110    0000010001001111    0000010001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01100 - 01104

  --0000010001010001    0000010001010010    0000010001010011    0000010001010100    0000010001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01105 - 01109

  --0000010001010110    0000010001010111    0000010001011000    0000010001011001    0000010001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01110 - 01114

  --0000010001011011    0000010001011100    0000010001011101    0000010001011110    0000010001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01115 - 01119

  --0000010001100000    0000010001100001    0000010001100010    0000010001100011    0000010001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01120 - 01124

  --0000010001100101    0000010001100110    0000010001100111    0000010001101000    0000010001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01125 - 01129

  --0000010001101010    0000010001101011    0000010001101100    0000010001101101    0000010001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01130 - 01134

  --0000010001101111    0000010001110000    0000010001110001    0000010001110010    0000010001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01135 - 01139

  --0000010001110100    0000010001110101    0000010001110110    0000010001110111    0000010001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01140 - 01144

  --0000010001111001    0000010001111010    0000010001111011    0000010001111100    0000010001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01145 - 01149

  --0000010001111110    0000010001111111    0000010010000000    0000010010000001    0000010010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01150 - 01154

  --0000010010000011    0000010010000100    0000010010000101    0000010010000110    0000010010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01155 - 01159

  --0000010010001000    0000010010001001    0000010010001010    0000010010001011    0000010010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01160 - 01164

  --0000010010001101    0000010010001110    0000010010001111    0000010010010000    0000010010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01165 - 01169

  --0000010010010010    0000010010010011    0000010010010100    0000010010010101    0000010010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01170 - 01174

  --0000010010010111    0000010010011000    0000010010011001    0000010010011010    0000010010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01175 - 01179

  --0000010010011100    0000010010011101    0000010010011110    0000010010011111    0000010010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01180 - 01184

  --0000010010100001    0000010010100010    0000010010100011    0000010010100100    0000010010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01185 - 01189

  --0000010010100110    0000010010100111    0000010010101000    0000010010101001    0000010010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01190 - 01194

  --0000010010101011    0000010010101100    0000010010101101    0000010010101110    0000010010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01195 - 01199

  --0000010010110000    0000010010110001    0000010010110010    0000010010110011    0000010010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01200 - 01204

  --0000010010110101    0000010010110110    0000010010110111    0000010010111000    0000010010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01205 - 01209

  --0000010010111010    0000010010111011    0000010010111100    0000010010111101    0000010010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01210 - 01214

  --0000010010111111    0000010011000000    0000010011000001    0000010011000010    0000010011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01215 - 01219

  --0000010011000100    0000010011000101    0000010011000110    0000010011000111    0000010011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01220 - 01224

  --0000010011001001    0000010011001010    0000010011001011    0000010011001100    0000010011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01225 - 01229

  --0000010011001110    0000010011001111    0000010011010000    0000010011010001    0000010011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01230 - 01234

  --0000010011010011    0000010011010100    0000010011010101    0000010011010110    0000010011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01235 - 01239

  --0000010011011000    0000010011011001    0000010011011010    0000010011011011    0000010011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01240 - 01244

  --0000010011011101    0000010011011110    0000010011011111    0000010011100000    0000010011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01245 - 01249

  --0000010011100010    0000010011100011    0000010011100100    0000010011100101    0000010011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01250 - 01254

  --0000010011100111    0000010011101000    0000010011101001    0000010011101010    0000010011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01255 - 01259

  --0000010011101100    0000010011101101    0000010011101110    0000010011101111    0000010011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01260 - 01264

  --0000010011110001    0000010011110010    0000010011110011    0000010011110100    0000010011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01265 - 01269

  --0000010011110110    0000010011110111    0000010011111000    0000010011111001    0000010011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01270 - 01274

  --0000010011111011    0000010011111100    0000010011111101    0000010011111110    0000010011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01275 - 01279

  --0000010100000000    0000010100000001    0000010100000010    0000010100000011    0000010100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01280 - 01284

  --0000010100000101    0000010100000110    0000010100000111    0000010100001000    0000010100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01285 - 01289

  --0000010100001010    0000010100001011    0000010100001100    0000010100001101    0000010100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01290 - 01294

  --0000010100001111    0000010100010000    0000010100010001    0000010100010010    0000010100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01295 - 01299

  --0000010100010100    0000010100010101    0000010100010110    0000010100010111    0000010100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01300 - 01304

  --0000010100011001    0000010100011010    0000010100011011    0000010100011100    0000010100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01305 - 01309

  --0000010100011110    0000010100011111    0000010100100000    0000010100100001    0000010100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01310 - 01314

  --0000010100100011    0000010100100100    0000010100100101    0000010100100110    0000010100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01315 - 01319

  --0000010100101000    0000010100101001    0000010100101010    0000010100101011    0000010100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01320 - 01324

  --0000010100101101    0000010100101110    0000010100101111    0000010100110000    0000010100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01325 - 01329

  --0000010100110010    0000010100110011    0000010100110100    0000010100110101    0000010100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01330 - 01334

  --0000010100110111    0000010100111000    0000010100111001    0000010100111010    0000010100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01335 - 01339

  --0000010100111100    0000010100111101    0000010100111110    0000010100111111    0000010101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01340 - 01344

  --0000010101000001    0000010101000010    0000010101000011    0000010101000100    0000010101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01345 - 01349

  --0000010101000110    0000010101000111    0000010101001000    0000010101001001    0000010101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01350 - 01354

  --0000010101001011    0000010101001100    0000010101001101    0000010101001110    0000010101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01355 - 01359

  --0000010101010000    0000010101010001    0000010101010010    0000010101010011    0000010101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01360 - 01364

  --0000010101010101    0000010101010110    0000010101010111    0000010101011000    0000010101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01365 - 01369

  --0000010101011010    0000010101011011    0000010101011100    0000010101011101    0000010101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01370 - 01374

  --0000010101011111    0000010101100000    0000010101100001    0000010101100010    0000010101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01375 - 01379

  --0000010101100100    0000010101100101    0000010101100110    0000010101100111    0000010101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01380 - 01384

  --0000010101101001    0000010101101010    0000010101101011    0000010101101100    0000010101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01385 - 01389

  --0000010101101110    0000010101101111    0000010101110000    0000010101110001    0000010101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01390 - 01394

  --0000010101110011    0000010101110100    0000010101110101    0000010101110110    0000010101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01395 - 01399

  --0000010101111000    0000010101111001    0000010101111010    0000010101111011    0000010101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01400 - 01404

  --0000010101111101    0000010101111110    0000010101111111    0000010110000000    0000010110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01405 - 01409

  --0000010110000010    0000010110000011    0000010110000100    0000010110000101    0000010110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01410 - 01414

  --0000010110000111    0000010110001000    0000010110001001    0000010110001010    0000010110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01415 - 01419

  --0000010110001100    0000010110001101    0000010110001110    0000010110001111    0000010110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01420 - 01424

  --0000010110010001    0000010110010010    0000010110010011    0000010110010100    0000010110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01425 - 01429

  --0000010110010110    0000010110010111    0000010110011000    0000010110011001    0000010110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01430 - 01434

  --0000010110011011    0000010110011100    0000010110011101    0000010110011110    0000010110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01435 - 01439

  --0000010110100000    0000010110100001    0000010110100010    0000010110100011    0000010110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01440 - 01444

  --0000010110100101    0000010110100110    0000010110100111    0000010110101000    0000010110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01445 - 01449

  --0000010110101010    0000010110101011    0000010110101100    0000010110101101    0000010110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01450 - 01454

  --0000010110101111    0000010110110000    0000010110110001    0000010110110010    0000010110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01455 - 01459

  --0000010110110100    0000010110110101    0000010110110110    0000010110110111    0000010110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01460 - 01464

  --0000010110111001    0000010110111010    0000010110111011    0000010110111100    0000010110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01465 - 01469

  --0000010110111110    0000010110111111    0000010111000000    0000010111000001    0000010111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01470 - 01474

  --0000010111000011    0000010111000100    0000010111000101    0000010111000110    0000010111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01475 - 01479

  --0000010111001000    0000010111001001    0000010111001010    0000010111001011    0000010111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01480 - 01484

  --0000010111001101    0000010111001110    0000010111001111    0000010111010000    0000010111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01485 - 01489

  --0000010111010010    0000010111010011    0000010111010100    0000010111010101    0000010111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01490 - 01494

  --0000010111010111    0000010111011000    0000010111011001    0000010111011010    0000010111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01495 - 01499

  --0000010111011100    0000010111011101    0000010111011110    0000010111011111    0000010111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01500 - 01504

  --0000010111100001    0000010111100010    0000010111100011    0000010111100100    0000010111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01505 - 01509

  --0000010111100110    0000010111100111    0000010111101000    0000010111101001    0000010111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01510 - 01514

  --0000010111101011    0000010111101100    0000010111101101    0000010111101110    0000010111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01515 - 01519

  --0000010111110000    0000010111110001    0000010111110010    0000010111110011    0000010111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01520 - 01524

  --0000010111110101    0000010111110110    0000010111110111    0000010111111000    0000010111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01525 - 01529

  --0000010111111010    0000010111111011    0000010111111100    0000010111111101    0000010111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01530 - 01534

  --0000010111111111    0000011000000000    0000011000000001    0000011000000010    0000011000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01535 - 01539

  --0000011000000100    0000011000000101    0000011000000110    0000011000000111    0000011000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01540 - 01544

  --0000011000001001    0000011000001010    0000011000001011    0000011000001100    0000011000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01545 - 01549

  --0000011000001110    0000011000001111    0000011000010000    0000011000010001    0000011000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01550 - 01554

  --0000011000010011    0000011000010100    0000011000010101    0000011000010110    0000011000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01555 - 01559

  --0000011000011000    0000011000011001    0000011000011010    0000011000011011    0000011000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01560 - 01564

  --0000011000011101    0000011000011110    0000011000011111    0000011000100000    0000011000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01565 - 01569

  --0000011000100010    0000011000100011    0000011000100100    0000011000100101    0000011000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01570 - 01574

  --0000011000100111    0000011000101000    0000011000101001    0000011000101010    0000011000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01575 - 01579

  --0000011000101100    0000011000101101    0000011000101110    0000011000101111    0000011000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01580 - 01584

  --0000011000110001    0000011000110010    0000011000110011    0000011000110100    0000011000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01585 - 01589

  --0000011000110110    0000011000110111    0000011000111000    0000011000111001    0000011000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01590 - 01594

  --0000011000111011    0000011000111100    0000011000111101    0000011000111110    0000011000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01595 - 01599

  --0000011001000000    0000011001000001    0000011001000010    0000011001000011    0000011001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01600 - 01604

  --0000011001000101    0000011001000110    0000011001000111    0000011001001000    0000011001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01605 - 01609

  --0000011001001010    0000011001001011    0000011001001100    0000011001001101    0000011001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01610 - 01614

  --0000011001001111    0000011001010000    0000011001010001    0000011001010010    0000011001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01615 - 01619

  --0000011001010100    0000011001010101    0000011001010110    0000011001010111    0000011001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01620 - 01624

  --0000011001011001    0000011001011010    0000011001011011    0000011001011100    0000011001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01625 - 01629

  --0000011001011110    0000011001011111    0000011001100000    0000011001100001    0000011001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01630 - 01634

  --0000011001100011    0000011001100100    0000011001100101    0000011001100110    0000011001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01635 - 01639

  --0000011001101000    0000011001101001    0000011001101010    0000011001101011    0000011001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01640 - 01644

  --0000011001101101    0000011001101110    0000011001101111    0000011001110000    0000011001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01645 - 01649

  --0000011001110010    0000011001110011    0000011001110100    0000011001110101    0000011001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01650 - 01654

  --0000011001110111    0000011001111000    0000011001111001    0000011001111010    0000011001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01655 - 01659

  --0000011001111100    0000011001111101    0000011001111110    0000011001111111    0000011010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01660 - 01664

  --0000011010000001    0000011010000010    0000011010000011    0000011010000100    0000011010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01665 - 01669

  --0000011010000110    0000011010000111    0000011010001000    0000011010001001    0000011010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01670 - 01674

  --0000011010001011    0000011010001100    0000011010001101    0000011010001110    0000011010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01675 - 01679

  --0000011010010000    0000011010010001    0000011010010010    0000011010010011    0000011010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01680 - 01684

  --0000011010010101    0000011010010110    0000011010010111    0000011010011000    0000011010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01685 - 01689

  --0000011010011010    0000011010011011    0000011010011100    0000011010011101    0000011010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01690 - 01694

  --0000011010011111    0000011010100000    0000011010100001    0000011010100010    0000011010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01695 - 01699

  --0000011010100100    0000011010100101    0000011010100110    0000011010100111    0000011010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01700 - 01704

  --0000011010101001    0000011010101010    0000011010101011    0000011010101100    0000011010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01705 - 01709

  --0000011010101110    0000011010101111    0000011010110000    0000011010110001    0000011010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01710 - 01714

  --0000011010110011    0000011010110100    0000011010110101    0000011010110110    0000011010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01715 - 01719

  --0000011010111000    0000011010111001    0000011010111010    0000011010111011    0000011010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01720 - 01724

  --0000011010111101    0000011010111110    0000011010111111    0000011011000000    0000011011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01725 - 01729

  --0000011011000010    0000011011000011    0000011011000100    0000011011000101    0000011011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01730 - 01734

  --0000011011000111    0000011011001000    0000011011001001    0000011011001010    0000011011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01735 - 01739

  --0000011011001100    0000011011001101    0000011011001110    0000011011001111    0000011011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01740 - 01744

  --0000011011010001    0000011011010010    0000011011010011    0000011011010100    0000011011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01745 - 01749

  --0000011011010110    0000011011010111    0000011011011000    0000011011011001    0000011011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01750 - 01754

  --0000011011011011    0000011011011100    0000011011011101    0000011011011110    0000011011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01755 - 01759

  --0000011011100000    0000011011100001    0000011011100010    0000011011100011    0000011011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01760 - 01764

  --0000011011100101    0000011011100110    0000011011100111    0000011011101000    0000011011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01765 - 01769

  --0000011011101010    0000011011101011    0000011011101100    0000011011101101    0000011011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01770 - 01774

  --0000011011101111    0000011011110000    0000011011110001    0000011011110010    0000011011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01775 - 01779

  --0000011011110100    0000011011110101    0000011011110110    0000011011110111    0000011011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01780 - 01784

  --0000011011111001    0000011011111010    0000011011111011    0000011011111100    0000011011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01785 - 01789

  --0000011011111110    0000011011111111    0000011100000000    0000011100000001    0000011100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01790 - 01794

  --0000011100000011    0000011100000100    0000011100000101    0000011100000110    0000011100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01795 - 01799

  --0000011100001000    0000011100001001    0000011100001010    0000011100001011    0000011100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01800 - 01804

  --0000011100001101    0000011100001110    0000011100001111    0000011100010000    0000011100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01805 - 01809

  --0000011100010010    0000011100010011    0000011100010100    0000011100010101    0000011100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01810 - 01814

  --0000011100010111    0000011100011000    0000011100011001    0000011100011010    0000011100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01815 - 01819

  --0000011100011100    0000011100011101    0000011100011110    0000011100011111    0000011100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01820 - 01824

  --0000011100100001    0000011100100010    0000011100100011    0000011100100100    0000011100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01825 - 01829

  --0000011100100110    0000011100100111    0000011100101000    0000011100101001    0000011100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01830 - 01834

  --0000011100101011    0000011100101100    0000011100101101    0000011100101110    0000011100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01835 - 01839

  --0000011100110000    0000011100110001    0000011100110010    0000011100110011    0000011100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01840 - 01844

  --0000011100110101    0000011100110110    0000011100110111    0000011100111000    0000011100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01845 - 01849

  --0000011100111010    0000011100111011    0000011100111100    0000011100111101    0000011100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01850 - 01854

  --0000011100111111    0000011101000000    0000011101000001    0000011101000010    0000011101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01855 - 01859

  --0000011101000100    0000011101000101    0000011101000110    0000011101000111    0000011101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01860 - 01864

  --0000011101001001    0000011101001010    0000011101001011    0000011101001100    0000011101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01865 - 01869

  --0000011101001110    0000011101001111    0000011101010000    0000011101010001    0000011101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01870 - 01874

  --0000011101010011    0000011101010100    0000011101010101    0000011101010110    0000011101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01875 - 01879

  --0000011101011000    0000011101011001    0000011101011010    0000011101011011    0000011101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01880 - 01884

  --0000011101011101    0000011101011110    0000011101011111    0000011101100000    0000011101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01885 - 01889

  --0000011101100010    0000011101100011    0000011101100100    0000011101100101    0000011101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01890 - 01894

  --0000011101100111    0000011101101000    0000011101101001    0000011101101010    0000011101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01895 - 01899

  --0000011101101100    0000011101101101    0000011101101110    0000011101101111    0000011101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01900 - 01904

  --0000011101110001    0000011101110010    0000011101110011    0000011101110100    0000011101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01905 - 01909

  --0000011101110110    0000011101110111    0000011101111000    0000011101111001    0000011101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01910 - 01914

  --0000011101111011    0000011101111100    0000011101111101    0000011101111110    0000011101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01915 - 01919

  --0000011110000000    0000011110000001    0000011110000010    0000011110000011    0000011110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01920 - 01924

  --0000011110000101    0000011110000110    0000011110000111    0000011110001000    0000011110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01925 - 01929

  --0000011110001010    0000011110001011    0000011110001100    0000011110001101    0000011110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01930 - 01934

  --0000011110001111    0000011110010000    0000011110010001    0000011110010010    0000011110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01935 - 01939

  --0000011110010100    0000011110010101    0000011110010110    0000011110010111    0000011110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01940 - 01944

  --0000011110011001    0000011110011010    0000011110011011    0000011110011100    0000011110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01945 - 01949

  --0000011110011110    0000011110011111    0000011110100000    0000011110100001    0000011110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01950 - 01954

  --0000011110100011    0000011110100100    0000011110100101    0000011110100110    0000011110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01955 - 01959

  --0000011110101000    0000011110101001    0000011110101010    0000011110101011    0000011110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01960 - 01964

  --0000011110101101    0000011110101110    0000011110101111    0000011110110000    0000011110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01965 - 01969

  --0000011110110010    0000011110110011    0000011110110100    0000011110110101    0000011110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01970 - 01974

  --0000011110110111    0000011110111000    0000011110111001    0000011110111010    0000011110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01975 - 01979

  --0000011110111100    0000011110111101    0000011110111110    0000011110111111    0000011111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01980 - 01984

  --0000011111000001    0000011111000010    0000011111000011    0000011111000100    0000011111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01985 - 01989

  --0000011111000110    0000011111000111    0000011111001000    0000011111001001    0000011111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01990 - 01994

  --0000011111001011    0000011111001100    0000011111001101    0000011111001110    0000011111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 01995 - 01999

  --0000011111010000    0000011111010001    0000011111010010    0000011111010011    0000011111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02000 - 02004

  --0000011111010101    0000011111010110    0000011111010111    0000011111011000    0000011111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02005 - 02009

  --0000011111011010    0000011111011011    0000011111011100    0000011111011101    0000011111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02010 - 02014

  --0000011111011111    0000011111100000    0000011111100001    0000011111100010    0000011111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02015 - 02019

  --0000011111100100    0000011111100101    0000011111100110    0000011111100111    0000011111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02020 - 02024

  --0000011111101001    0000011111101010    0000011111101011    0000011111101100    0000011111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02025 - 02029

  --0000011111101110    0000011111101111    0000011111110000    0000011111110001    0000011111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02030 - 02034

  --0000011111110011    0000011111110100    0000011111110101    0000011111110110    0000011111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02035 - 02039

  --0000011111111000    0000011111111001    0000011111111010    0000011111111011    0000011111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02040 - 02044

  --0000011111111101    0000011111111110    0000011111111111    0000100000000000    0000100000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02045 - 02049

  --0000100000000010    0000100000000011    0000100000000100    0000100000000101    0000100000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02050 - 02054

  --0000100000000111    0000100000001000    0000100000001001    0000100000001010    0000100000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02055 - 02059

  --0000100000001100    0000100000001101    0000100000001110    0000100000001111    0000100000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02060 - 02064

  --0000100000010001    0000100000010010    0000100000010011    0000100000010100    0000100000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02065 - 02069

  --0000100000010110    0000100000010111    0000100000011000    0000100000011001    0000100000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02070 - 02074

  --0000100000011011    0000100000011100    0000100000011101    0000100000011110    0000100000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02075 - 02079

  --0000100000100000    0000100000100001    0000100000100010    0000100000100011    0000100000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02080 - 02084

  --0000100000100101    0000100000100110    0000100000100111    0000100000101000    0000100000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02085 - 02089

  --0000100000101010    0000100000101011    0000100000101100    0000100000101101    0000100000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02090 - 02094

  --0000100000101111    0000100000110000    0000100000110001    0000100000110010    0000100000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02095 - 02099

  --0000100000110100    0000100000110101    0000100000110110    0000100000110111    0000100000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02100 - 02104

  --0000100000111001    0000100000111010    0000100000111011    0000100000111100    0000100000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02105 - 02109

  --0000100000111110    0000100000111111    0000100001000000    0000100001000001    0000100001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02110 - 02114

  --0000100001000011    0000100001000100    0000100001000101    0000100001000110    0000100001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02115 - 02119

  --0000100001001000    0000100001001001    0000100001001010    0000100001001011    0000100001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02120 - 02124

  --0000100001001101    0000100001001110    0000100001001111    0000100001010000    0000100001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02125 - 02129

  --0000100001010010    0000100001010011    0000100001010100    0000100001010101    0000100001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02130 - 02134

  --0000100001010111    0000100001011000    0000100001011001    0000100001011010    0000100001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02135 - 02139

  --0000100001011100    0000100001011101    0000100001011110    0000100001011111    0000100001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02140 - 02144

  --0000100001100001    0000100001100010    0000100001100011    0000100001100100    0000100001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02145 - 02149

  --0000100001100110    0000100001100111    0000100001101000    0000100001101001    0000100001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02150 - 02154

  --0000100001101011    0000100001101100    0000100001101101    0000100001101110    0000100001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02155 - 02159

  --0000100001110000    0000100001110001    0000100001110010    0000100001110011    0000100001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02160 - 02164

  --0000100001110101    0000100001110110    0000100001110111    0000100001111000    0000100001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02165 - 02169

  --0000100001111010    0000100001111011    0000100001111100    0000100001111101    0000100001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02170 - 02174

  --0000100001111111    0000100010000000    0000100010000001    0000100010000010    0000100010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02175 - 02179

  --0000100010000100    0000100010000101    0000100010000110    0000100010000111    0000100010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02180 - 02184

  --0000100010001001    0000100010001010    0000100010001011    0000100010001100    0000100010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02185 - 02189

  --0000100010001110    0000100010001111    0000100010010000    0000100010010001    0000100010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02190 - 02194

  --0000100010010011    0000100010010100    0000100010010101    0000100010010110    0000100010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02195 - 02199

  --0000100010011000    0000100010011001    0000100010011010    0000100010011011    0000100010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02200 - 02204

  --0000100010011101    0000100010011110    0000100010011111    0000100010100000    0000100010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02205 - 02209

  --0000100010100010    0000100010100011    0000100010100100    0000100010100101    0000100010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02210 - 02214

  --0000100010100111    0000100010101000    0000100010101001    0000100010101010    0000100010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02215 - 02219

  --0000100010101100    0000100010101101    0000100010101110    0000100010101111    0000100010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02220 - 02224

  --0000100010110001    0000100010110010    0000100010110011    0000100010110100    0000100010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02225 - 02229

  --0000100010110110    0000100010110111    0000100010111000    0000100010111001    0000100010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02230 - 02234

  --0000100010111011    0000100010111100    0000100010111101    0000100010111110    0000100010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02235 - 02239

  --0000100011000000    0000100011000001    0000100011000010    0000100011000011    0000100011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02240 - 02244

  --0000100011000101    0000100011000110    0000100011000111    0000100011001000    0000100011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02245 - 02249

  --0000100011001010    0000100011001011    0000100011001100    0000100011001101    0000100011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02250 - 02254

  --0000100011001111    0000100011010000    0000100011010001    0000100011010010    0000100011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02255 - 02259

  --0000100011010100    0000100011010101    0000100011010110    0000100011010111    0000100011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02260 - 02264

  --0000100011011001    0000100011011010    0000100011011011    0000100011011100    0000100011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02265 - 02269

  --0000100011011110    0000100011011111    0000100011100000    0000100011100001    0000100011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02270 - 02274

  --0000100011100011    0000100011100100    0000100011100101    0000100011100110    0000100011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02275 - 02279

  --0000100011101000    0000100011101001    0000100011101010    0000100011101011    0000100011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02280 - 02284

  --0000100011101101    0000100011101110    0000100011101111    0000100011110000    0000100011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02285 - 02289

  --0000100011110010    0000100011110011    0000100011110100    0000100011110101    0000100011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02290 - 02294

  --0000100011110111    0000100011111000    0000100011111001    0000100011111010    0000100011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02295 - 02299

  --0000100011111100    0000100011111101    0000100011111110    0000100011111111    0000100100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02300 - 02304

  --0000100100000001    0000100100000010    0000100100000011    0000100100000100    0000100100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02305 - 02309

  --0000100100000110    0000100100000111    0000100100001000    0000100100001001    0000100100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02310 - 02314

  --0000100100001011    0000100100001100    0000100100001101    0000100100001110    0000100100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02315 - 02319

  --0000100100010000    0000100100010001    0000100100010010    0000100100010011    0000100100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02320 - 02324

  --0000100100010101    0000100100010110    0000100100010111    0000100100011000    0000100100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02325 - 02329

  --0000100100011010    0000100100011011    0000100100011100    0000100100011101    0000100100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02330 - 02334

  --0000100100011111    0000100100100000    0000100100100001    0000100100100010    0000100100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02335 - 02339

  --0000100100100100    0000100100100101    0000100100100110    0000100100100111    0000100100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02340 - 02344

  --0000100100101001    0000100100101010    0000100100101011    0000100100101100    0000100100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02345 - 02349

  --0000100100101110    0000100100101111    0000100100110000    0000100100110001    0000100100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02350 - 02354

  --0000100100110011    0000100100110100    0000100100110101    0000100100110110    0000100100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02355 - 02359

  --0000100100111000    0000100100111001    0000100100111010    0000100100111011    0000100100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02360 - 02364

  --0000100100111101    0000100100111110    0000100100111111    0000100101000000    0000100101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02365 - 02369

  --0000100101000010    0000100101000011    0000100101000100    0000100101000101    0000100101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02370 - 02374

  --0000100101000111    0000100101001000    0000100101001001    0000100101001010    0000100101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02375 - 02379

  --0000100101001100    0000100101001101    0000100101001110    0000100101001111    0000100101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02380 - 02384

  --0000100101010001    0000100101010010    0000100101010011    0000100101010100    0000100101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02385 - 02389

  --0000100101010110    0000100101010111    0000100101011000    0000100101011001    0000100101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02390 - 02394

  --0000100101011011    0000100101011100    0000100101011101    0000100101011110    0000100101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02395 - 02399

  --0000100101100000    0000100101100001    0000100101100010    0000100101100011    0000100101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02400 - 02404

  --0000100101100101    0000100101100110    0000100101100111    0000100101101000    0000100101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02405 - 02409

  --0000100101101010    0000100101101011    0000100101101100    0000100101101101    0000100101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02410 - 02414

  --0000100101101111    0000100101110000    0000100101110001    0000100101110010    0000100101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02415 - 02419

  --0000100101110100    0000100101110101    0000100101110110    0000100101110111    0000100101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02420 - 02424

  --0000100101111001    0000100101111010    0000100101111011    0000100101111100    0000100101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02425 - 02429

  --0000100101111110    0000100101111111    0000100110000000    0000100110000001    0000100110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02430 - 02434

  --0000100110000011    0000100110000100    0000100110000101    0000100110000110    0000100110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02435 - 02439

  --0000100110001000    0000100110001001    0000100110001010    0000100110001011    0000100110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02440 - 02444

  --0000100110001101    0000100110001110    0000100110001111    0000100110010000    0000100110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02445 - 02449

  --0000100110010010    0000100110010011    0000100110010100    0000100110010101    0000100110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02450 - 02454

  --0000100110010111    0000100110011000    0000100110011001    0000100110011010    0000100110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02455 - 02459

  --0000100110011100    0000100110011101    0000100110011110    0000100110011111    0000100110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02460 - 02464

  --0000100110100001    0000100110100010    0000100110100011    0000100110100100    0000100110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02465 - 02469

  --0000100110100110    0000100110100111    0000100110101000    0000100110101001    0000100110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02470 - 02474

  --0000100110101011    0000100110101100    0000100110101101    0000100110101110    0000100110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02475 - 02479

  --0000100110110000    0000100110110001    0000100110110010    0000100110110011    0000100110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02480 - 02484

  --0000100110110101    0000100110110110    0000100110110111    0000100110111000    0000100110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02485 - 02489

  --0000100110111010    0000100110111011    0000100110111100    0000100110111101    0000100110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02490 - 02494

  --0000100110111111    0000100111000000    0000100111000001    0000100111000010    0000100111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02495 - 02499

  --0000100111000100    0000100111000101    0000100111000110    0000100111000111    0000100111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02500 - 02504

  --0000100111001001    0000100111001010    0000100111001011    0000100111001100    0000100111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02505 - 02509

  --0000100111001110    0000100111001111    0000100111010000    0000100111010001    0000100111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02510 - 02514

  --0000100111010011    0000100111010100    0000100111010101    0000100111010110    0000100111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02515 - 02519

  --0000100111011000    0000100111011001    0000100111011010    0000100111011011    0000100111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02520 - 02524

  --0000100111011101    0000100111011110    0000100111011111    0000100111100000    0000100111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02525 - 02529

  --0000100111100010    0000100111100011    0000100111100100    0000100111100101    0000100111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02530 - 02534

  --0000100111100111    0000100111101000    0000100111101001    0000100111101010    0000100111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02535 - 02539

  --0000100111101100    0000100111101101    0000100111101110    0000100111101111    0000100111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02540 - 02544

  --0000100111110001    0000100111110010    0000100111110011    0000100111110100    0000100111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02545 - 02549

  --0000100111110110    0000100111110111    0000100111111000    0000100111111001    0000100111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02550 - 02554

  --0000100111111011    0000100111111100    0000100111111101    0000100111111110    0000100111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02555 - 02559

  --0000101000000000    0000101000000001    0000101000000010    0000101000000011    0000101000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02560 - 02564

  --0000101000000101    0000101000000110    0000101000000111    0000101000001000    0000101000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02565 - 02569

  --0000101000001010    0000101000001011    0000101000001100    0000101000001101    0000101000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02570 - 02574

  --0000101000001111    0000101000010000    0000101000010001    0000101000010010    0000101000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02575 - 02579

  --0000101000010100    0000101000010101    0000101000010110    0000101000010111    0000101000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02580 - 02584

  --0000101000011001    0000101000011010    0000101000011011    0000101000011100    0000101000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02585 - 02589

  --0000101000011110    0000101000011111    0000101000100000    0000101000100001    0000101000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02590 - 02594

  --0000101000100011    0000101000100100    0000101000100101    0000101000100110    0000101000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02595 - 02599

  --0000101000101000    0000101000101001    0000101000101010    0000101000101011    0000101000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02600 - 02604

  --0000101000101101    0000101000101110    0000101000101111    0000101000110000    0000101000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02605 - 02609

  --0000101000110010    0000101000110011    0000101000110100    0000101000110101    0000101000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02610 - 02614

  --0000101000110111    0000101000111000    0000101000111001    0000101000111010    0000101000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02615 - 02619

  --0000101000111100    0000101000111101    0000101000111110    0000101000111111    0000101001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02620 - 02624

  --0000101001000001    0000101001000010    0000101001000011    0000101001000100    0000101001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02625 - 02629

  --0000101001000110    0000101001000111    0000101001001000    0000101001001001    0000101001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02630 - 02634

  --0000101001001011    0000101001001100    0000101001001101    0000101001001110    0000101001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02635 - 02639

  --0000101001010000    0000101001010001    0000101001010010    0000101001010011    0000101001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02640 - 02644

  --0000101001010101    0000101001010110    0000101001010111    0000101001011000    0000101001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02645 - 02649

  --0000101001011010    0000101001011011    0000101001011100    0000101001011101    0000101001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02650 - 02654

  --0000101001011111    0000101001100000    0000101001100001    0000101001100010    0000101001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02655 - 02659

  --0000101001100100    0000101001100101    0000101001100110    0000101001100111    0000101001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02660 - 02664

  --0000101001101001    0000101001101010    0000101001101011    0000101001101100    0000101001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02665 - 02669

  --0000101001101110    0000101001101111    0000101001110000    0000101001110001    0000101001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02670 - 02674

  --0000101001110011    0000101001110100    0000101001110101    0000101001110110    0000101001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02675 - 02679

  --0000101001111000    0000101001111001    0000101001111010    0000101001111011    0000101001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02680 - 02684

  --0000101001111101    0000101001111110    0000101001111111    0000101010000000    0000101010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02685 - 02689

  --0000101010000010    0000101010000011    0000101010000100    0000101010000101    0000101010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02690 - 02694

  --0000101010000111    0000101010001000    0000101010001001    0000101010001010    0000101010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02695 - 02699

  --0000101010001100    0000101010001101    0000101010001110    0000101010001111    0000101010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02700 - 02704

  --0000101010010001    0000101010010010    0000101010010011    0000101010010100    0000101010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02705 - 02709

  --0000101010010110    0000101010010111    0000101010011000    0000101010011001    0000101010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02710 - 02714

  --0000101010011011    0000101010011100    0000101010011101    0000101010011110    0000101010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02715 - 02719

  --0000101010100000    0000101010100001    0000101010100010    0000101010100011    0000101010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02720 - 02724

  --0000101010100101    0000101010100110    0000101010100111    0000101010101000    0000101010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02725 - 02729

  --0000101010101010    0000101010101011    0000101010101100    0000101010101101    0000101010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02730 - 02734

  --0000101010101111    0000101010110000    0000101010110001    0000101010110010    0000101010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02735 - 02739

  --0000101010110100    0000101010110101    0000101010110110    0000101010110111    0000101010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02740 - 02744

  --0000101010111001    0000101010111010    0000101010111011    0000101010111100    0000101010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02745 - 02749

  --0000101010111110    0000101010111111    0000101011000000    0000101011000001    0000101011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02750 - 02754

  --0000101011000011    0000101011000100    0000101011000101    0000101011000110    0000101011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02755 - 02759

  --0000101011001000    0000101011001001    0000101011001010    0000101011001011    0000101011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02760 - 02764

  --0000101011001101    0000101011001110    0000101011001111    0000101011010000    0000101011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02765 - 02769

  --0000101011010010    0000101011010011    0000101011010100    0000101011010101    0000101011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02770 - 02774

  --0000101011010111    0000101011011000    0000101011011001    0000101011011010    0000101011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02775 - 02779

  --0000101011011100    0000101011011101    0000101011011110    0000101011011111    0000101011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02780 - 02784

  --0000101011100001    0000101011100010    0000101011100011    0000101011100100    0000101011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02785 - 02789

  --0000101011100110    0000101011100111    0000101011101000    0000101011101001    0000101011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02790 - 02794

  --0000101011101011    0000101011101100    0000101011101101    0000101011101110    0000101011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02795 - 02799

  --0000101011110000    0000101011110001    0000101011110010    0000101011110011    0000101011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02800 - 02804

  --0000101011110101    0000101011110110    0000101011110111    0000101011111000    0000101011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02805 - 02809

  --0000101011111010    0000101011111011    0000101011111100    0000101011111101    0000101011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02810 - 02814

  --0000101011111111    0000101100000000    0000101100000001    0000101100000010    0000101100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02815 - 02819

  --0000101100000100    0000101100000101    0000101100000110    0000101100000111    0000101100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02820 - 02824

  --0000101100001001    0000101100001010    0000101100001011    0000101100001100    0000101100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02825 - 02829

  --0000101100001110    0000101100001111    0000101100010000    0000101100010001    0000101100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02830 - 02834

  --0000101100010011    0000101100010100    0000101100010101    0000101100010110    0000101100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02835 - 02839

  --0000101100011000    0000101100011001    0000101100011010    0000101100011011    0000101100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02840 - 02844

  --0000101100011101    0000101100011110    0000101100011111    0000101100100000    0000101100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02845 - 02849

  --0000101100100010    0000101100100011    0000101100100100    0000101100100101    0000101100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02850 - 02854

  --0000101100100111    0000101100101000    0000101100101001    0000101100101010    0000101100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02855 - 02859

  --0000101100101100    0000101100101101    0000101100101110    0000101100101111    0000101100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02860 - 02864

  --0000101100110001    0000101100110010    0000101100110011    0000101100110100    0000101100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02865 - 02869

  --0000101100110110    0000101100110111    0000101100111000    0000101100111001    0000101100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02870 - 02874

  --0000101100111011    0000101100111100    0000101100111101    0000101100111110    0000101100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02875 - 02879

  --0000101101000000    0000101101000001    0000101101000010    0000101101000011    0000101101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02880 - 02884

  --0000101101000101    0000101101000110    0000101101000111    0000101101001000    0000101101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02885 - 02889

  --0000101101001010    0000101101001011    0000101101001100    0000101101001101    0000101101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02890 - 02894

  --0000101101001111    0000101101010000    0000101101010001    0000101101010010    0000101101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02895 - 02899

  --0000101101010100    0000101101010101    0000101101010110    0000101101010111    0000101101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02900 - 02904

  --0000101101011001    0000101101011010    0000101101011011    0000101101011100    0000101101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02905 - 02909

  --0000101101011110    0000101101011111    0000101101100000    0000101101100001    0000101101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02910 - 02914

  --0000101101100011    0000101101100100    0000101101100101    0000101101100110    0000101101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02915 - 02919

  --0000101101101000    0000101101101001    0000101101101010    0000101101101011    0000101101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02920 - 02924

  --0000101101101101    0000101101101110    0000101101101111    0000101101110000    0000101101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02925 - 02929

  --0000101101110010    0000101101110011    0000101101110100    0000101101110101    0000101101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02930 - 02934

  --0000101101110111    0000101101111000    0000101101111001    0000101101111010    0000101101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02935 - 02939

  --0000101101111100    0000101101111101    0000101101111110    0000101101111111    0000101110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02940 - 02944

  --0000101110000001    0000101110000010    0000101110000011    0000101110000100    0000101110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02945 - 02949

  --0000101110000110    0000101110000111    0000101110001000    0000101110001001    0000101110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02950 - 02954

  --0000101110001011    0000101110001100    0000101110001101    0000101110001110    0000101110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02955 - 02959

  --0000101110010000    0000101110010001    0000101110010010    0000101110010011    0000101110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02960 - 02964

  --0000101110010101    0000101110010110    0000101110010111    0000101110011000    0000101110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02965 - 02969

  --0000101110011010    0000101110011011    0000101110011100    0000101110011101    0000101110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02970 - 02974

  --0000101110011111    0000101110100000    0000101110100001    0000101110100010    0000101110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02975 - 02979

  --0000101110100100    0000101110100101    0000101110100110    0000101110100111    0000101110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02980 - 02984

  --0000101110101001    0000101110101010    0000101110101011    0000101110101100    0000101110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02985 - 02989

  --0000101110101110    0000101110101111    0000101110110000    0000101110110001    0000101110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02990 - 02994

  --0000101110110011    0000101110110100    0000101110110101    0000101110110110    0000101110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 02995 - 02999

  --0000101110111000    0000101110111001    0000101110111010    0000101110111011    0000101110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03000 - 03004

  --0000101110111101    0000101110111110    0000101110111111    0000101111000000    0000101111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03005 - 03009

  --0000101111000010    0000101111000011    0000101111000100    0000101111000101    0000101111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03010 - 03014

  --0000101111000111    0000101111001000    0000101111001001    0000101111001010    0000101111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03015 - 03019

  --0000101111001100    0000101111001101    0000101111001110    0000101111001111    0000101111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03020 - 03024

  --0000101111010001    0000101111010010    0000101111010011    0000101111010100    0000101111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03025 - 03029

  --0000101111010110    0000101111010111    0000101111011000    0000101111011001    0000101111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03030 - 03034

  --0000101111011011    0000101111011100    0000101111011101    0000101111011110    0000101111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03035 - 03039

  --0000101111100000    0000101111100001    0000101111100010    0000101111100011    0000101111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03040 - 03044

  --0000101111100101    0000101111100110    0000101111100111    0000101111101000    0000101111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03045 - 03049

  --0000101111101010    0000101111101011    0000101111101100    0000101111101101    0000101111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03050 - 03054

  --0000101111101111    0000101111110000    0000101111110001    0000101111110010    0000101111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03055 - 03059

  --0000101111110100    0000101111110101    0000101111110110    0000101111110111    0000101111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03060 - 03064

  --0000101111111001    0000101111111010    0000101111111011    0000101111111100    0000101111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03065 - 03069

  --0000101111111110    0000101111111111    0000110000000000    0000110000000001    0000110000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03070 - 03074

  --0000110000000011    0000110000000100    0000110000000101    0000110000000110    0000110000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03075 - 03079

  --0000110000001000    0000110000001001    0000110000001010    0000110000001011    0000110000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03080 - 03084

  --0000110000001101    0000110000001110    0000110000001111    0000110000010000    0000110000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03085 - 03089

  --0000110000010010    0000110000010011    0000110000010100    0000110000010101    0000110000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03090 - 03094

  --0000110000010111    0000110000011000    0000110000011001    0000110000011010    0000110000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03095 - 03099

  --0000110000011100    0000110000011101    0000110000011110    0000110000011111    0000110000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03100 - 03104

  --0000110000100001    0000110000100010    0000110000100011    0000110000100100    0000110000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03105 - 03109

  --0000110000100110    0000110000100111    0000110000101000    0000110000101001    0000110000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03110 - 03114

  --0000110000101011    0000110000101100    0000110000101101    0000110000101110    0000110000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03115 - 03119

  --0000110000110000    0000110000110001    0000110000110010    0000110000110011    0000110000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03120 - 03124

  --0000110000110101    0000110000110110    0000110000110111    0000110000111000    0000110000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03125 - 03129

  --0000110000111010    0000110000111011    0000110000111100    0000110000111101    0000110000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03130 - 03134

  --0000110000111111    0000110001000000    0000110001000001    0000110001000010    0000110001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03135 - 03139

  --0000110001000100    0000110001000101    0000110001000110    0000110001000111    0000110001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03140 - 03144

  --0000110001001001    0000110001001010    0000110001001011    0000110001001100    0000110001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03145 - 03149

  --0000110001001110    0000110001001111    0000110001010000    0000110001010001    0000110001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03150 - 03154

  --0000110001010011    0000110001010100    0000110001010101    0000110001010110    0000110001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03155 - 03159

  --0000110001011000    0000110001011001    0000110001011010    0000110001011011    0000110001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03160 - 03164

  --0000110001011101    0000110001011110    0000110001011111    0000110001100000    0000110001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03165 - 03169

  --0000110001100010    0000110001100011    0000110001100100    0000110001100101    0000110001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03170 - 03174

  --0000110001100111    0000110001101000    0000110001101001    0000110001101010    0000110001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03175 - 03179

  --0000110001101100    0000110001101101    0000110001101110    0000110001101111    0000110001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03180 - 03184

  --0000110001110001    0000110001110010    0000110001110011    0000110001110100    0000110001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03185 - 03189

  --0000110001110110    0000110001110111    0000110001111000    0000110001111001    0000110001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03190 - 03194

  --0000110001111011    0000110001111100    0000110001111101    0000110001111110    0000110001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03195 - 03199

  --0000110010000000    0000110010000001    0000110010000010    0000110010000011    0000110010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03200 - 03204

  --0000110010000101    0000110010000110    0000110010000111    0000110010001000    0000110010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03205 - 03209

  --0000110010001010    0000110010001011    0000110010001100    0000110010001101    0000110010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03210 - 03214

  --0000110010001111    0000110010010000    0000110010010001    0000110010010010    0000110010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03215 - 03219

  --0000110010010100    0000110010010101    0000110010010110    0000110010010111    0000110010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03220 - 03224

  --0000110010011001    0000110010011010    0000110010011011    0000110010011100    0000110010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03225 - 03229

  --0000110010011110    0000110010011111    0000110010100000    0000110010100001    0000110010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03230 - 03234

  --0000110010100011    0000110010100100    0000110010100101    0000110010100110    0000110010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03235 - 03239

  --0000110010101000    0000110010101001    0000110010101010    0000110010101011    0000110010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03240 - 03244

  --0000110010101101    0000110010101110    0000110010101111    0000110010110000    0000110010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03245 - 03249

  --0000110010110010    0000110010110011    0000110010110100    0000110010110101    0000110010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03250 - 03254

  --0000110010110111    0000110010111000    0000110010111001    0000110010111010    0000110010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03255 - 03259

  --0000110010111100    0000110010111101    0000110010111110    0000110010111111    0000110011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03260 - 03264

  --0000110011000001    0000110011000010    0000110011000011    0000110011000100    0000110011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03265 - 03269

  --0000110011000110    0000110011000111    0000110011001000    0000110011001001    0000110011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03270 - 03274

  --0000110011001011    0000110011001100    0000110011001101    0000110011001110    0000110011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03275 - 03279

  --0000110011010000    0000110011010001    0000110011010010    0000110011010011    0000110011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03280 - 03284

  --0000110011010101    0000110011010110    0000110011010111    0000110011011000    0000110011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03285 - 03289

  --0000110011011010    0000110011011011    0000110011011100    0000110011011101    0000110011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03290 - 03294

  --0000110011011111    0000110011100000    0000110011100001    0000110011100010    0000110011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03295 - 03299

  --0000110011100100    0000110011100101    0000110011100110    0000110011100111    0000110011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03300 - 03304

  --0000110011101001    0000110011101010    0000110011101011    0000110011101100    0000110011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03305 - 03309

  --0000110011101110    0000110011101111    0000110011110000    0000110011110001    0000110011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03310 - 03314

  --0000110011110011    0000110011110100    0000110011110101    0000110011110110    0000110011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03315 - 03319

  --0000110011111000    0000110011111001    0000110011111010    0000110011111011    0000110011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03320 - 03324

  --0000110011111101    0000110011111110    0000110011111111    0000110100000000    0000110100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03325 - 03329

  --0000110100000010    0000110100000011    0000110100000100    0000110100000101    0000110100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03330 - 03334

  --0000110100000111    0000110100001000    0000110100001001    0000110100001010    0000110100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03335 - 03339

  --0000110100001100    0000110100001101    0000110100001110    0000110100001111    0000110100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03340 - 03344

  --0000110100010001    0000110100010010    0000110100010011    0000110100010100    0000110100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03345 - 03349

  --0000110100010110    0000110100010111    0000110100011000    0000110100011001    0000110100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03350 - 03354

  --0000110100011011    0000110100011100    0000110100011101    0000110100011110    0000110100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03355 - 03359

  --0000110100100000    0000110100100001    0000110100100010    0000110100100011    0000110100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03360 - 03364

  --0000110100100101    0000110100100110    0000110100100111    0000110100101000    0000110100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03365 - 03369

  --0000110100101010    0000110100101011    0000110100101100    0000110100101101    0000110100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03370 - 03374

  --0000110100101111    0000110100110000    0000110100110001    0000110100110010    0000110100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03375 - 03379

  --0000110100110100    0000110100110101    0000110100110110    0000110100110111    0000110100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03380 - 03384

  --0000110100111001    0000110100111010    0000110100111011    0000110100111100    0000110100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03385 - 03389

  --0000110100111110    0000110100111111    0000110101000000    0000110101000001    0000110101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03390 - 03394

  --0000110101000011    0000110101000100    0000110101000101    0000110101000110    0000110101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03395 - 03399

  --0000110101001000    0000110101001001    0000110101001010    0000110101001011    0000110101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03400 - 03404

  --0000110101001101    0000110101001110    0000110101001111    0000110101010000    0000110101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03405 - 03409

  --0000110101010010    0000110101010011    0000110101010100    0000110101010101    0000110101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03410 - 03414

  --0000110101010111    0000110101011000    0000110101011001    0000110101011010    0000110101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03415 - 03419

  --0000110101011100    0000110101011101    0000110101011110    0000110101011111    0000110101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03420 - 03424

  --0000110101100001    0000110101100010    0000110101100011    0000110101100100    0000110101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03425 - 03429

  --0000110101100110    0000110101100111    0000110101101000    0000110101101001    0000110101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03430 - 03434

  --0000110101101011    0000110101101100    0000110101101101    0000110101101110    0000110101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03435 - 03439

  --0000110101110000    0000110101110001    0000110101110010    0000110101110011    0000110101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03440 - 03444

  --0000110101110101    0000110101110110    0000110101110111    0000110101111000    0000110101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03445 - 03449

  --0000110101111010    0000110101111011    0000110101111100    0000110101111101    0000110101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03450 - 03454

  --0000110101111111    0000110110000000    0000110110000001    0000110110000010    0000110110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03455 - 03459

  --0000110110000100    0000110110000101    0000110110000110    0000110110000111    0000110110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03460 - 03464

  --0000110110001001    0000110110001010    0000110110001011    0000110110001100    0000110110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03465 - 03469

  --0000110110001110    0000110110001111    0000110110010000    0000110110010001    0000110110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03470 - 03474

  --0000110110010011    0000110110010100    0000110110010101    0000110110010110    0000110110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03475 - 03479

  --0000110110011000    0000110110011001    0000110110011010    0000110110011011    0000110110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03480 - 03484

  --0000110110011101    0000110110011110    0000110110011111    0000110110100000    0000110110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03485 - 03489

  --0000110110100010    0000110110100011    0000110110100100    0000110110100101    0000110110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03490 - 03494

  --0000110110100111    0000110110101000    0000110110101001    0000110110101010    0000110110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03495 - 03499

  --0000110110101100    0000110110101101    0000110110101110    0000110110101111    0000110110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03500 - 03504

  --0000110110110001    0000110110110010    0000110110110011    0000110110110100    0000110110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03505 - 03509

  --0000110110110110    0000110110110111    0000110110111000    0000110110111001    0000110110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03510 - 03514

  --0000110110111011    0000110110111100    0000110110111101    0000110110111110    0000110110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03515 - 03519

  --0000110111000000    0000110111000001    0000110111000010    0000110111000011    0000110111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03520 - 03524

  --0000110111000101    0000110111000110    0000110111000111    0000110111001000    0000110111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03525 - 03529

  --0000110111001010    0000110111001011    0000110111001100    0000110111001101    0000110111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03530 - 03534

  --0000110111001111    0000110111010000    0000110111010001    0000110111010010    0000110111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03535 - 03539

  --0000110111010100    0000110111010101    0000110111010110    0000110111010111    0000110111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03540 - 03544

  --0000110111011001    0000110111011010    0000110111011011    0000110111011100    0000110111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03545 - 03549

  --0000110111011110    0000110111011111    0000110111100000    0000110111100001    0000110111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03550 - 03554

  --0000110111100011    0000110111100100    0000110111100101    0000110111100110    0000110111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03555 - 03559

  --0000110111101000    0000110111101001    0000110111101010    0000110111101011    0000110111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03560 - 03564

  --0000110111101101    0000110111101110    0000110111101111    0000110111110000    0000110111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03565 - 03569

  --0000110111110010    0000110111110011    0000110111110100    0000110111110101    0000110111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03570 - 03574

  --0000110111110111    0000110111111000    0000110111111001    0000110111111010    0000110111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03575 - 03579

  --0000110111111100    0000110111111101    0000110111111110    0000110111111111    0000111000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03580 - 03584

  --0000111000000001    0000111000000010    0000111000000011    0000111000000100    0000111000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03585 - 03589

  --0000111000000110    0000111000000111    0000111000001000    0000111000001001    0000111000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03590 - 03594

  --0000111000001011    0000111000001100    0000111000001101    0000111000001110    0000111000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03595 - 03599

  --0000111000010000    0000111000010001    0000111000010010    0000111000010011    0000111000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03600 - 03604

  --0000111000010101    0000111000010110    0000111000010111    0000111000011000    0000111000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03605 - 03609

  --0000111000011010    0000111000011011    0000111000011100    0000111000011101    0000111000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03610 - 03614

  --0000111000011111    0000111000100000    0000111000100001    0000111000100010    0000111000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03615 - 03619

  --0000111000100100    0000111000100101    0000111000100110    0000111000100111    0000111000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03620 - 03624

  --0000111000101001    0000111000101010    0000111000101011    0000111000101100    0000111000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03625 - 03629

  --0000111000101110    0000111000101111    0000111000110000    0000111000110001    0000111000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03630 - 03634

  --0000111000110011    0000111000110100    0000111000110101    0000111000110110    0000111000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03635 - 03639

  --0000111000111000    0000111000111001    0000111000111010    0000111000111011    0000111000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03640 - 03644

  --0000111000111101    0000111000111110    0000111000111111    0000111001000000    0000111001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03645 - 03649

  --0000111001000010    0000111001000011    0000111001000100    0000111001000101    0000111001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03650 - 03654

  --0000111001000111    0000111001001000    0000111001001001    0000111001001010    0000111001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03655 - 03659

  --0000111001001100    0000111001001101    0000111001001110    0000111001001111    0000111001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03660 - 03664

  --0000111001010001    0000111001010010    0000111001010011    0000111001010100    0000111001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03665 - 03669

  --0000111001010110    0000111001010111    0000111001011000    0000111001011001    0000111001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03670 - 03674

  --0000111001011011    0000111001011100    0000111001011101    0000111001011110    0000111001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03675 - 03679

  --0000111001100000    0000111001100001    0000111001100010    0000111001100011    0000111001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03680 - 03684

  --0000111001100101    0000111001100110    0000111001100111    0000111001101000    0000111001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03685 - 03689

  --0000111001101010    0000111001101011    0000111001101100    0000111001101101    0000111001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03690 - 03694

  --0000111001101111    0000111001110000    0000111001110001    0000111001110010    0000111001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03695 - 03699

  --0000111001110100    0000111001110101    0000111001110110    0000111001110111    0000111001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03700 - 03704

  --0000111001111001    0000111001111010    0000111001111011    0000111001111100    0000111001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03705 - 03709

  --0000111001111110    0000111001111111    0000111010000000    0000111010000001    0000111010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03710 - 03714

  --0000111010000011    0000111010000100    0000111010000101    0000111010000110    0000111010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03715 - 03719

  --0000111010001000    0000111010001001    0000111010001010    0000111010001011    0000111010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03720 - 03724

  --0000111010001101    0000111010001110    0000111010001111    0000111010010000    0000111010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03725 - 03729

  --0000111010010010    0000111010010011    0000111010010100    0000111010010101    0000111010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03730 - 03734

  --0000111010010111    0000111010011000    0000111010011001    0000111010011010    0000111010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03735 - 03739

  --0000111010011100    0000111010011101    0000111010011110    0000111010011111    0000111010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03740 - 03744

  --0000111010100001    0000111010100010    0000111010100011    0000111010100100    0000111010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03745 - 03749

  --0000111010100110    0000111010100111    0000111010101000    0000111010101001    0000111010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03750 - 03754

  --0000111010101011    0000111010101100    0000111010101101    0000111010101110    0000111010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03755 - 03759

  --0000111010110000    0000111010110001    0000111010110010    0000111010110011    0000111010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03760 - 03764

  --0000111010110101    0000111010110110    0000111010110111    0000111010111000    0000111010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03765 - 03769

  --0000111010111010    0000111010111011    0000111010111100    0000111010111101    0000111010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03770 - 03774

  --0000111010111111    0000111011000000    0000111011000001    0000111011000010    0000111011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03775 - 03779

  --0000111011000100    0000111011000101    0000111011000110    0000111011000111    0000111011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03780 - 03784

  --0000111011001001    0000111011001010    0000111011001011    0000111011001100    0000111011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03785 - 03789

  --0000111011001110    0000111011001111    0000111011010000    0000111011010001    0000111011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03790 - 03794

  --0000111011010011    0000111011010100    0000111011010101    0000111011010110    0000111011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03795 - 03799

  --0000111011011000    0000111011011001    0000111011011010    0000111011011011    0000111011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03800 - 03804

  --0000111011011101    0000111011011110    0000111011011111    0000111011100000    0000111011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03805 - 03809

  --0000111011100010    0000111011100011    0000111011100100    0000111011100101    0000111011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03810 - 03814

  --0000111011100111    0000111011101000    0000111011101001    0000111011101010    0000111011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03815 - 03819

  --0000111011101100    0000111011101101    0000111011101110    0000111011101111    0000111011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03820 - 03824

  --0000111011110001    0000111011110010    0000111011110011    0000111011110100    0000111011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03825 - 03829

  --0000111011110110    0000111011110111    0000111011111000    0000111011111001    0000111011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03830 - 03834

  --0000111011111011    0000111011111100    0000111011111101    0000111011111110    0000111011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03835 - 03839

  --0000111100000000    0000111100000001    0000111100000010    0000111100000011    0000111100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03840 - 03844

  --0000111100000101    0000111100000110    0000111100000111    0000111100001000    0000111100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03845 - 03849

  --0000111100001010    0000111100001011    0000111100001100    0000111100001101    0000111100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03850 - 03854

  --0000111100001111    0000111100010000    0000111100010001    0000111100010010    0000111100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03855 - 03859

  --0000111100010100    0000111100010101    0000111100010110    0000111100010111    0000111100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03860 - 03864

  --0000111100011001    0000111100011010    0000111100011011    0000111100011100    0000111100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03865 - 03869

  --0000111100011110    0000111100011111    0000111100100000    0000111100100001    0000111100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03870 - 03874

  --0000111100100011    0000111100100100    0000111100100101    0000111100100110    0000111100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03875 - 03879

  --0000111100101000    0000111100101001    0000111100101010    0000111100101011    0000111100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03880 - 03884

  --0000111100101101    0000111100101110    0000111100101111    0000111100110000    0000111100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03885 - 03889

  --0000111100110010    0000111100110011    0000111100110100    0000111100110101    0000111100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03890 - 03894

  --0000111100110111    0000111100111000    0000111100111001    0000111100111010    0000111100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03895 - 03899

  --0000111100111100    0000111100111101    0000111100111110    0000111100111111    0000111101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03900 - 03904

  --0000111101000001    0000111101000010    0000111101000011    0000111101000100    0000111101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03905 - 03909

  --0000111101000110    0000111101000111    0000111101001000    0000111101001001    0000111101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03910 - 03914

  --0000111101001011    0000111101001100    0000111101001101    0000111101001110    0000111101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03915 - 03919

  --0000111101010000    0000111101010001    0000111101010010    0000111101010011    0000111101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03920 - 03924

  --0000111101010101    0000111101010110    0000111101010111    0000111101011000    0000111101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03925 - 03929

  --0000111101011010    0000111101011011    0000111101011100    0000111101011101    0000111101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03930 - 03934

  --0000111101011111    0000111101100000    0000111101100001    0000111101100010    0000111101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03935 - 03939

  --0000111101100100    0000111101100101    0000111101100110    0000111101100111    0000111101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03940 - 03944

  --0000111101101001    0000111101101010    0000111101101011    0000111101101100    0000111101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03945 - 03949

  --0000111101101110    0000111101101111    0000111101110000    0000111101110001    0000111101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03950 - 03954

  --0000111101110011    0000111101110100    0000111101110101    0000111101110110    0000111101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03955 - 03959

  --0000111101111000    0000111101111001    0000111101111010    0000111101111011    0000111101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03960 - 03964

  --0000111101111101    0000111101111110    0000111101111111    0000111110000000    0000111110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03965 - 03969

  --0000111110000010    0000111110000011    0000111110000100    0000111110000101    0000111110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03970 - 03974

  --0000111110000111    0000111110001000    0000111110001001    0000111110001010    0000111110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03975 - 03979

  --0000111110001100    0000111110001101    0000111110001110    0000111110001111    0000111110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03980 - 03984

  --0000111110010001    0000111110010010    0000111110010011    0000111110010100    0000111110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03985 - 03989

  --0000111110010110    0000111110010111    0000111110011000    0000111110011001    0000111110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03990 - 03994

  --0000111110011011    0000111110011100    0000111110011101    0000111110011110    0000111110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 03995 - 03999

  --0000111110100000    0000111110100001    0000111110100010    0000111110100011    0000111110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04000 - 04004

  --0000111110100101    0000111110100110    0000111110100111    0000111110101000    0000111110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04005 - 04009

  --0000111110101010    0000111110101011    0000111110101100    0000111110101101    0000111110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04010 - 04014

  --0000111110101111    0000111110110000    0000111110110001    0000111110110010    0000111110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04015 - 04019

  --0000111110110100    0000111110110101    0000111110110110    0000111110110111    0000111110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04020 - 04024

  --0000111110111001    0000111110111010    0000111110111011    0000111110111100    0000111110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04025 - 04029

  --0000111110111110    0000111110111111    0000111111000000    0000111111000001    0000111111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04030 - 04034

  --0000111111000011    0000111111000100    0000111111000101    0000111111000110    0000111111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04035 - 04039

  --0000111111001000    0000111111001001    0000111111001010    0000111111001011    0000111111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04040 - 04044

  --0000111111001101    0000111111001110    0000111111001111    0000111111010000    0000111111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04045 - 04049

  --0000111111010010    0000111111010011    0000111111010100    0000111111010101    0000111111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04050 - 04054

  --0000111111010111    0000111111011000    0000111111011001    0000111111011010    0000111111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04055 - 04059

  --0000111111011100    0000111111011101    0000111111011110    0000111111011111    0000111111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04060 - 04064

  --0000111111100001    0000111111100010    0000111111100011    0000111111100100    0000111111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04065 - 04069

  --0000111111100110    0000111111100111    0000111111101000    0000111111101001    0000111111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04070 - 04074

  --0000111111101011    0000111111101100    0000111111101101    0000111111101110    0000111111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04075 - 04079

  --0000111111110000    0000111111110001    0000111111110010    0000111111110011    0000111111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04080 - 04084

  --0000111111110101    0000111111110110    0000111111110111    0000111111111000    0000111111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04085 - 04089

  --0000111111111010    0000111111111011    0000111111111100    0000111111111101    0000111111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04090 - 04094

  --0000111111111111    0001000000000000    0001000000000001    0001000000000010    0001000000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04095 - 04099

  --0001000000000100    0001000000000101    0001000000000110    0001000000000111    0001000000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04100 - 04104

  --0001000000001001    0001000000001010    0001000000001011    0001000000001100    0001000000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04105 - 04109

  --0001000000001110    0001000000001111    0001000000010000    0001000000010001    0001000000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04110 - 04114

  --0001000000010011    0001000000010100    0001000000010101    0001000000010110    0001000000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04115 - 04119

  --0001000000011000    0001000000011001    0001000000011010    0001000000011011    0001000000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04120 - 04124

  --0001000000011101    0001000000011110    0001000000011111    0001000000100000    0001000000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04125 - 04129

  --0001000000100010    0001000000100011    0001000000100100    0001000000100101    0001000000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04130 - 04134

  --0001000000100111    0001000000101000    0001000000101001    0001000000101010    0001000000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04135 - 04139

  --0001000000101100    0001000000101101    0001000000101110    0001000000101111    0001000000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04140 - 04144

  --0001000000110001    0001000000110010    0001000000110011    0001000000110100    0001000000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04145 - 04149

  --0001000000110110    0001000000110111    0001000000111000    0001000000111001    0001000000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04150 - 04154

  --0001000000111011    0001000000111100    0001000000111101    0001000000111110    0001000000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04155 - 04159

  --0001000001000000    0001000001000001    0001000001000010    0001000001000011    0001000001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04160 - 04164

  --0001000001000101    0001000001000110    0001000001000111    0001000001001000    0001000001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04165 - 04169

  --0001000001001010    0001000001001011    0001000001001100    0001000001001101    0001000001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04170 - 04174

  --0001000001001111    0001000001010000    0001000001010001    0001000001010010    0001000001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04175 - 04179

  --0001000001010100    0001000001010101    0001000001010110    0001000001010111    0001000001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04180 - 04184

  --0001000001011001    0001000001011010    0001000001011011    0001000001011100    0001000001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04185 - 04189

  --0001000001011110    0001000001011111    0001000001100000    0001000001100001    0001000001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04190 - 04194

  --0001000001100011    0001000001100100    0001000001100101    0001000001100110    0001000001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04195 - 04199

  --0001000001101000    0001000001101001    0001000001101010    0001000001101011    0001000001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04200 - 04204

  --0001000001101101    0001000001101110    0001000001101111    0001000001110000    0001000001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04205 - 04209

  --0001000001110010    0001000001110011    0001000001110100    0001000001110101    0001000001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04210 - 04214

  --0001000001110111    0001000001111000    0001000001111001    0001000001111010    0001000001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04215 - 04219

  --0001000001111100    0001000001111101    0001000001111110    0001000001111111    0001000010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04220 - 04224

  --0001000010000001    0001000010000010    0001000010000011    0001000010000100    0001000010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04225 - 04229

  --0001000010000110    0001000010000111    0001000010001000    0001000010001001    0001000010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04230 - 04234

  --0001000010001011    0001000010001100    0001000010001101    0001000010001110    0001000010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04235 - 04239

  --0001000010010000    0001000010010001    0001000010010010    0001000010010011    0001000010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04240 - 04244

  --0001000010010101    0001000010010110    0001000010010111    0001000010011000    0001000010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04245 - 04249

  --0001000010011010    0001000010011011    0001000010011100    0001000010011101    0001000010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04250 - 04254

  --0001000010011111    0001000010100000    0001000010100001    0001000010100010    0001000010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04255 - 04259

  --0001000010100100    0001000010100101    0001000010100110    0001000010100111    0001000010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04260 - 04264

  --0001000010101001    0001000010101010    0001000010101011    0001000010101100    0001000010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04265 - 04269

  --0001000010101110    0001000010101111    0001000010110000    0001000010110001    0001000010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04270 - 04274

  --0001000010110011    0001000010110100    0001000010110101    0001000010110110    0001000010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04275 - 04279

  --0001000010111000    0001000010111001    0001000010111010    0001000010111011    0001000010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04280 - 04284

  --0001000010111101    0001000010111110    0001000010111111    0001000011000000    0001000011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04285 - 04289

  --0001000011000010    0001000011000011    0001000011000100    0001000011000101    0001000011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04290 - 04294

  --0001000011000111    0001000011001000    0001000011001001    0001000011001010    0001000011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04295 - 04299

  --0001000011001100    0001000011001101    0001000011001110    0001000011001111    0001000011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04300 - 04304

  --0001000011010001    0001000011010010    0001000011010011    0001000011010100    0001000011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04305 - 04309

  --0001000011010110    0001000011010111    0001000011011000    0001000011011001    0001000011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04310 - 04314

  --0001000011011011    0001000011011100    0001000011011101    0001000011011110    0001000011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04315 - 04319

  --0001000011100000    0001000011100001    0001000011100010    0001000011100011    0001000011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04320 - 04324

  --0001000011100101    0001000011100110    0001000011100111    0001000011101000    0001000011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04325 - 04329

  --0001000011101010    0001000011101011    0001000011101100    0001000011101101    0001000011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04330 - 04334

  --0001000011101111    0001000011110000    0001000011110001    0001000011110010    0001000011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04335 - 04339

  --0001000011110100    0001000011110101    0001000011110110    0001000011110111    0001000011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04340 - 04344

  --0001000011111001    0001000011111010    0001000011111011    0001000011111100    0001000011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04345 - 04349

  --0001000011111110    0001000011111111    0001000100000000    0001000100000001    0001000100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04350 - 04354

  --0001000100000011    0001000100000100    0001000100000101    0001000100000110    0001000100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04355 - 04359

  --0001000100001000    0001000100001001    0001000100001010    0001000100001011    0001000100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04360 - 04364

  --0001000100001101    0001000100001110    0001000100001111    0001000100010000    0001000100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04365 - 04369

  --0001000100010010    0001000100010011    0001000100010100    0001000100010101    0001000100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04370 - 04374

  --0001000100010111    0001000100011000    0001000100011001    0001000100011010    0001000100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04375 - 04379

  --0001000100011100    0001000100011101    0001000100011110    0001000100011111    0001000100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04380 - 04384

  --0001000100100001    0001000100100010    0001000100100011    0001000100100100    0001000100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04385 - 04389

  --0001000100100110    0001000100100111    0001000100101000    0001000100101001    0001000100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04390 - 04394

  --0001000100101011    0001000100101100    0001000100101101    0001000100101110    0001000100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04395 - 04399

  --0001000100110000    0001000100110001    0001000100110010    0001000100110011    0001000100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04400 - 04404

  --0001000100110101    0001000100110110    0001000100110111    0001000100111000    0001000100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04405 - 04409

  --0001000100111010    0001000100111011    0001000100111100    0001000100111101    0001000100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04410 - 04414

  --0001000100111111    0001000101000000    0001000101000001    0001000101000010    0001000101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04415 - 04419

  --0001000101000100    0001000101000101    0001000101000110    0001000101000111    0001000101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04420 - 04424

  --0001000101001001    0001000101001010    0001000101001011    0001000101001100    0001000101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04425 - 04429

  --0001000101001110    0001000101001111    0001000101010000    0001000101010001    0001000101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04430 - 04434

  --0001000101010011    0001000101010100    0001000101010101    0001000101010110    0001000101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04435 - 04439

  --0001000101011000    0001000101011001    0001000101011010    0001000101011011    0001000101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04440 - 04444

  --0001000101011101    0001000101011110    0001000101011111    0001000101100000    0001000101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04445 - 04449

  --0001000101100010    0001000101100011    0001000101100100    0001000101100101    0001000101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04450 - 04454

  --0001000101100111    0001000101101000    0001000101101001    0001000101101010    0001000101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04455 - 04459

  --0001000101101100    0001000101101101    0001000101101110    0001000101101111    0001000101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04460 - 04464

  --0001000101110001    0001000101110010    0001000101110011    0001000101110100    0001000101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04465 - 04469

  --0001000101110110    0001000101110111    0001000101111000    0001000101111001    0001000101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04470 - 04474

  --0001000101111011    0001000101111100    0001000101111101    0001000101111110    0001000101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04475 - 04479

  --0001000110000000    0001000110000001    0001000110000010    0001000110000011    0001000110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04480 - 04484

  --0001000110000101    0001000110000110    0001000110000111    0001000110001000    0001000110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04485 - 04489

  --0001000110001010    0001000110001011    0001000110001100    0001000110001101    0001000110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04490 - 04494

  --0001000110001111    0001000110010000    0001000110010001    0001000110010010    0001000110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04495 - 04499

  --0001000110010100    0001000110010101    0001000110010110    0001000110010111    0001000110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04500 - 04504

  --0001000110011001    0001000110011010    0001000110011011    0001000110011100    0001000110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04505 - 04509

  --0001000110011110    0001000110011111    0001000110100000    0001000110100001    0001000110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04510 - 04514

  --0001000110100011    0001000110100100    0001000110100101    0001000110100110    0001000110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04515 - 04519

  --0001000110101000    0001000110101001    0001000110101010    0001000110101011    0001000110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04520 - 04524

  --0001000110101101    0001000110101110    0001000110101111    0001000110110000    0001000110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04525 - 04529

  --0001000110110010    0001000110110011    0001000110110100    0001000110110101    0001000110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04530 - 04534

  --0001000110110111    0001000110111000    0001000110111001    0001000110111010    0001000110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04535 - 04539

  --0001000110111100    0001000110111101    0001000110111110    0001000110111111    0001000111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04540 - 04544

  --0001000111000001    0001000111000010    0001000111000011    0001000111000100    0001000111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04545 - 04549

  --0001000111000110    0001000111000111    0001000111001000    0001000111001001    0001000111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04550 - 04554

  --0001000111001011    0001000111001100    0001000111001101    0001000111001110    0001000111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04555 - 04559

  --0001000111010000    0001000111010001    0001000111010010    0001000111010011    0001000111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04560 - 04564

  --0001000111010101    0001000111010110    0001000111010111    0001000111011000    0001000111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04565 - 04569

  --0001000111011010    0001000111011011    0001000111011100    0001000111011101    0001000111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04570 - 04574

  --0001000111011111    0001000111100000    0001000111100001    0001000111100010    0001000111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04575 - 04579

  --0001000111100100    0001000111100101    0001000111100110    0001000111100111    0001000111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04580 - 04584

  --0001000111101001    0001000111101010    0001000111101011    0001000111101100    0001000111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04585 - 04589

  --0001000111101110    0001000111101111    0001000111110000    0001000111110001    0001000111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04590 - 04594

  --0001000111110011    0001000111110100    0001000111110101    0001000111110110    0001000111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04595 - 04599

  --0001000111111000    0001000111111001    0001000111111010    0001000111111011    0001000111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04600 - 04604

  --0001000111111101    0001000111111110    0001000111111111    0001001000000000    0001001000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04605 - 04609

  --0001001000000010    0001001000000011    0001001000000100    0001001000000101    0001001000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04610 - 04614

  --0001001000000111    0001001000001000    0001001000001001    0001001000001010    0001001000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04615 - 04619

  --0001001000001100    0001001000001101    0001001000001110    0001001000001111    0001001000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04620 - 04624

  --0001001000010001    0001001000010010    0001001000010011    0001001000010100    0001001000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04625 - 04629

  --0001001000010110    0001001000010111    0001001000011000    0001001000011001    0001001000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04630 - 04634

  --0001001000011011    0001001000011100    0001001000011101    0001001000011110    0001001000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04635 - 04639

  --0001001000100000    0001001000100001    0001001000100010    0001001000100011    0001001000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04640 - 04644

  --0001001000100101    0001001000100110    0001001000100111    0001001000101000    0001001000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04645 - 04649

  --0001001000101010    0001001000101011    0001001000101100    0001001000101101    0001001000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04650 - 04654

  --0001001000101111    0001001000110000    0001001000110001    0001001000110010    0001001000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04655 - 04659

  --0001001000110100    0001001000110101    0001001000110110    0001001000110111    0001001000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04660 - 04664

  --0001001000111001    0001001000111010    0001001000111011    0001001000111100    0001001000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04665 - 04669

  --0001001000111110    0001001000111111    0001001001000000    0001001001000001    0001001001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04670 - 04674

  --0001001001000011    0001001001000100    0001001001000101    0001001001000110    0001001001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04675 - 04679

  --0001001001001000    0001001001001001    0001001001001010    0001001001001011    0001001001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04680 - 04684

  --0001001001001101    0001001001001110    0001001001001111    0001001001010000    0001001001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04685 - 04689

  --0001001001010010    0001001001010011    0001001001010100    0001001001010101    0001001001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04690 - 04694

  --0001001001010111    0001001001011000    0001001001011001    0001001001011010    0001001001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04695 - 04699

  --0001001001011100    0001001001011101    0001001001011110    0001001001011111    0001001001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04700 - 04704

  --0001001001100001    0001001001100010    0001001001100011    0001001001100100    0001001001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04705 - 04709

  --0001001001100110    0001001001100111    0001001001101000    0001001001101001    0001001001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04710 - 04714

  --0001001001101011    0001001001101100    0001001001101101    0001001001101110    0001001001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04715 - 04719

  --0001001001110000    0001001001110001    0001001001110010    0001001001110011    0001001001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04720 - 04724

  --0001001001110101    0001001001110110    0001001001110111    0001001001111000    0001001001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04725 - 04729

  --0001001001111010    0001001001111011    0001001001111100    0001001001111101    0001001001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04730 - 04734

  --0001001001111111    0001001010000000    0001001010000001    0001001010000010    0001001010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04735 - 04739

  --0001001010000100    0001001010000101    0001001010000110    0001001010000111    0001001010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04740 - 04744

  --0001001010001001    0001001010001010    0001001010001011    0001001010001100    0001001010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04745 - 04749

  --0001001010001110    0001001010001111    0001001010010000    0001001010010001    0001001010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04750 - 04754

  --0001001010010011    0001001010010100    0001001010010101    0001001010010110    0001001010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04755 - 04759

  --0001001010011000    0001001010011001    0001001010011010    0001001010011011    0001001010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04760 - 04764

  --0001001010011101    0001001010011110    0001001010011111    0001001010100000    0001001010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04765 - 04769

  --0001001010100010    0001001010100011    0001001010100100    0001001010100101    0001001010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04770 - 04774

  --0001001010100111    0001001010101000    0001001010101001    0001001010101010    0001001010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04775 - 04779

  --0001001010101100    0001001010101101    0001001010101110    0001001010101111    0001001010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04780 - 04784

  --0001001010110001    0001001010110010    0001001010110011    0001001010110100    0001001010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04785 - 04789

  --0001001010110110    0001001010110111    0001001010111000    0001001010111001    0001001010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04790 - 04794

  --0001001010111011    0001001010111100    0001001010111101    0001001010111110    0001001010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04795 - 04799

  --0001001011000000    0001001011000001    0001001011000010    0001001011000011    0001001011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04800 - 04804

  --0001001011000101    0001001011000110    0001001011000111    0001001011001000    0001001011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04805 - 04809

  --0001001011001010    0001001011001011    0001001011001100    0001001011001101    0001001011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04810 - 04814

  --0001001011001111    0001001011010000    0001001011010001    0001001011010010    0001001011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04815 - 04819

  --0001001011010100    0001001011010101    0001001011010110    0001001011010111    0001001011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04820 - 04824

  --0001001011011001    0001001011011010    0001001011011011    0001001011011100    0001001011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04825 - 04829

  --0001001011011110    0001001011011111    0001001011100000    0001001011100001    0001001011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04830 - 04834

  --0001001011100011    0001001011100100    0001001011100101    0001001011100110    0001001011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04835 - 04839

  --0001001011101000    0001001011101001    0001001011101010    0001001011101011    0001001011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04840 - 04844

  --0001001011101101    0001001011101110    0001001011101111    0001001011110000    0001001011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04845 - 04849

  --0001001011110010    0001001011110011    0001001011110100    0001001011110101    0001001011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04850 - 04854

  --0001001011110111    0001001011111000    0001001011111001    0001001011111010    0001001011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04855 - 04859

  --0001001011111100    0001001011111101    0001001011111110    0001001011111111    0001001100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04860 - 04864

  --0001001100000001    0001001100000010    0001001100000011    0001001100000100    0001001100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04865 - 04869

  --0001001100000110    0001001100000111    0001001100001000    0001001100001001    0001001100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04870 - 04874

  --0001001100001011    0001001100001100    0001001100001101    0001001100001110    0001001100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04875 - 04879

  --0001001100010000    0001001100010001    0001001100010010    0001001100010011    0001001100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04880 - 04884

  --0001001100010101    0001001100010110    0001001100010111    0001001100011000    0001001100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04885 - 04889

  --0001001100011010    0001001100011011    0001001100011100    0001001100011101    0001001100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04890 - 04894

  --0001001100011111    0001001100100000    0001001100100001    0001001100100010    0001001100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04895 - 04899

  --0001001100100100    0001001100100101    0001001100100110    0001001100100111    0001001100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04900 - 04904

  --0001001100101001    0001001100101010    0001001100101011    0001001100101100    0001001100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04905 - 04909

  --0001001100101110    0001001100101111    0001001100110000    0001001100110001    0001001100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04910 - 04914

  --0001001100110011    0001001100110100    0001001100110101    0001001100110110    0001001100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04915 - 04919

  --0001001100111000    0001001100111001    0001001100111010    0001001100111011    0001001100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04920 - 04924

  --0001001100111101    0001001100111110    0001001100111111    0001001101000000    0001001101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04925 - 04929

  --0001001101000010    0001001101000011    0001001101000100    0001001101000101    0001001101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04930 - 04934

  --0001001101000111    0001001101001000    0001001101001001    0001001101001010    0001001101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04935 - 04939

  --0001001101001100    0001001101001101    0001001101001110    0001001101001111    0001001101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04940 - 04944

  --0001001101010001    0001001101010010    0001001101010011    0001001101010100    0001001101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04945 - 04949

  --0001001101010110    0001001101010111    0001001101011000    0001001101011001    0001001101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04950 - 04954

  --0001001101011011    0001001101011100    0001001101011101    0001001101011110    0001001101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04955 - 04959

  --0001001101100000    0001001101100001    0001001101100010    0001001101100011    0001001101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04960 - 04964

  --0001001101100101    0001001101100110    0001001101100111    0001001101101000    0001001101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04965 - 04969

  --0001001101101010    0001001101101011    0001001101101100    0001001101101101    0001001101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04970 - 04974

  --0001001101101111    0001001101110000    0001001101110001    0001001101110010    0001001101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04975 - 04979

  --0001001101110100    0001001101110101    0001001101110110    0001001101110111    0001001101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04980 - 04984

  --0001001101111001    0001001101111010    0001001101111011    0001001101111100    0001001101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04985 - 04989

  --0001001101111110    0001001101111111    0001001110000000    0001001110000001    0001001110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04990 - 04994

  --0001001110000011    0001001110000100    0001001110000101    0001001110000110    0001001110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 04995 - 04999

  --0001001110001000    0001001110001001    0001001110001010    0001001110001011    0001001110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05000 - 05004

  --0001001110001101    0001001110001110    0001001110001111    0001001110010000    0001001110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05005 - 05009

  --0001001110010010    0001001110010011    0001001110010100    0001001110010101    0001001110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05010 - 05014

  --0001001110010111    0001001110011000    0001001110011001    0001001110011010    0001001110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05015 - 05019

  --0001001110011100    0001001110011101    0001001110011110    0001001110011111    0001001110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05020 - 05024

  --0001001110100001    0001001110100010    0001001110100011    0001001110100100    0001001110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05025 - 05029

  --0001001110100110    0001001110100111    0001001110101000    0001001110101001    0001001110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05030 - 05034

  --0001001110101011    0001001110101100    0001001110101101    0001001110101110    0001001110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05035 - 05039

  --0001001110110000    0001001110110001    0001001110110010    0001001110110011    0001001110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05040 - 05044

  --0001001110110101    0001001110110110    0001001110110111    0001001110111000    0001001110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05045 - 05049

  --0001001110111010    0001001110111011    0001001110111100    0001001110111101    0001001110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05050 - 05054

  --0001001110111111    0001001111000000    0001001111000001    0001001111000010    0001001111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05055 - 05059

  --0001001111000100    0001001111000101    0001001111000110    0001001111000111    0001001111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05060 - 05064

  --0001001111001001    0001001111001010    0001001111001011    0001001111001100    0001001111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05065 - 05069

  --0001001111001110    0001001111001111    0001001111010000    0001001111010001    0001001111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05070 - 05074

  --0001001111010011    0001001111010100    0001001111010101    0001001111010110    0001001111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05075 - 05079

  --0001001111011000    0001001111011001    0001001111011010    0001001111011011    0001001111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05080 - 05084

  --0001001111011101    0001001111011110    0001001111011111    0001001111100000    0001001111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05085 - 05089

  --0001001111100010    0001001111100011    0001001111100100    0001001111100101    0001001111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05090 - 05094

  --0001001111100111    0001001111101000    0001001111101001    0001001111101010    0001001111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05095 - 05099

  --0001001111101100    0001001111101101    0001001111101110    0001001111101111    0001001111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05100 - 05104

  --0001001111110001    0001001111110010    0001001111110011    0001001111110100    0001001111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05105 - 05109

  --0001001111110110    0001001111110111    0001001111111000    0001001111111001    0001001111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05110 - 05114

  --0001001111111011    0001001111111100    0001001111111101    0001001111111110    0001001111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05115 - 05119

  --0001010000000000    0001010000000001    0001010000000010    0001010000000011    0001010000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05120 - 05124

  --0001010000000101    0001010000000110    0001010000000111    0001010000001000    0001010000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05125 - 05129

  --0001010000001010    0001010000001011    0001010000001100    0001010000001101    0001010000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05130 - 05134

  --0001010000001111    0001010000010000    0001010000010001    0001010000010010    0001010000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05135 - 05139

  --0001010000010100    0001010000010101    0001010000010110    0001010000010111    0001010000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05140 - 05144

  --0001010000011001    0001010000011010    0001010000011011    0001010000011100    0001010000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05145 - 05149

  --0001010000011110    0001010000011111    0001010000100000    0001010000100001    0001010000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05150 - 05154

  --0001010000100011    0001010000100100    0001010000100101    0001010000100110    0001010000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05155 - 05159

  --0001010000101000    0001010000101001    0001010000101010    0001010000101011    0001010000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05160 - 05164

  --0001010000101101    0001010000101110    0001010000101111    0001010000110000    0001010000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05165 - 05169

  --0001010000110010    0001010000110011    0001010000110100    0001010000110101    0001010000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05170 - 05174

  --0001010000110111    0001010000111000    0001010000111001    0001010000111010    0001010000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05175 - 05179

  --0001010000111100    0001010000111101    0001010000111110    0001010000111111    0001010001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05180 - 05184

  --0001010001000001    0001010001000010    0001010001000011    0001010001000100    0001010001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05185 - 05189

  --0001010001000110    0001010001000111    0001010001001000    0001010001001001    0001010001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05190 - 05194

  --0001010001001011    0001010001001100    0001010001001101    0001010001001110    0001010001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05195 - 05199

  --0001010001010000    0001010001010001    0001010001010010    0001010001010011    0001010001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05200 - 05204

  --0001010001010101    0001010001010110    0001010001010111    0001010001011000    0001010001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05205 - 05209

  --0001010001011010    0001010001011011    0001010001011100    0001010001011101    0001010001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05210 - 05214

  --0001010001011111    0001010001100000    0001010001100001    0001010001100010    0001010001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05215 - 05219

  --0001010001100100    0001010001100101    0001010001100110    0001010001100111    0001010001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05220 - 05224

  --0001010001101001    0001010001101010    0001010001101011    0001010001101100    0001010001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05225 - 05229

  --0001010001101110    0001010001101111    0001010001110000    0001010001110001    0001010001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05230 - 05234

  --0001010001110011    0001010001110100    0001010001110101    0001010001110110    0001010001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05235 - 05239

  --0001010001111000    0001010001111001    0001010001111010    0001010001111011    0001010001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05240 - 05244

  --0001010001111101    0001010001111110    0001010001111111    0001010010000000    0001010010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05245 - 05249

  --0001010010000010    0001010010000011    0001010010000100    0001010010000101    0001010010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05250 - 05254

  --0001010010000111    0001010010001000    0001010010001001    0001010010001010    0001010010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05255 - 05259

  --0001010010001100    0001010010001101    0001010010001110    0001010010001111    0001010010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05260 - 05264

  --0001010010010001    0001010010010010    0001010010010011    0001010010010100    0001010010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05265 - 05269

  --0001010010010110    0001010010010111    0001010010011000    0001010010011001    0001010010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05270 - 05274

  --0001010010011011    0001010010011100    0001010010011101    0001010010011110    0001010010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05275 - 05279

  --0001010010100000    0001010010100001    0001010010100010    0001010010100011    0001010010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05280 - 05284

  --0001010010100101    0001010010100110    0001010010100111    0001010010101000    0001010010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05285 - 05289

  --0001010010101010    0001010010101011    0001010010101100    0001010010101101    0001010010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05290 - 05294

  --0001010010101111    0001010010110000    0001010010110001    0001010010110010    0001010010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05295 - 05299

  --0001010010110100    0001010010110101    0001010010110110    0001010010110111    0001010010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05300 - 05304

  --0001010010111001    0001010010111010    0001010010111011    0001010010111100    0001010010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05305 - 05309

  --0001010010111110    0001010010111111    0001010011000000    0001010011000001    0001010011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05310 - 05314

  --0001010011000011    0001010011000100    0001010011000101    0001010011000110    0001010011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05315 - 05319

  --0001010011001000    0001010011001001    0001010011001010    0001010011001011    0001010011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05320 - 05324

  --0001010011001101    0001010011001110    0001010011001111    0001010011010000    0001010011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05325 - 05329

  --0001010011010010    0001010011010011    0001010011010100    0001010011010101    0001010011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05330 - 05334

  --0001010011010111    0001010011011000    0001010011011001    0001010011011010    0001010011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05335 - 05339

  --0001010011011100    0001010011011101    0001010011011110    0001010011011111    0001010011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05340 - 05344

  --0001010011100001    0001010011100010    0001010011100011    0001010011100100    0001010011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05345 - 05349

  --0001010011100110    0001010011100111    0001010011101000    0001010011101001    0001010011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05350 - 05354

  --0001010011101011    0001010011101100    0001010011101101    0001010011101110    0001010011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05355 - 05359

  --0001010011110000    0001010011110001    0001010011110010    0001010011110011    0001010011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05360 - 05364

  --0001010011110101    0001010011110110    0001010011110111    0001010011111000    0001010011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05365 - 05369

  --0001010011111010    0001010011111011    0001010011111100    0001010011111101    0001010011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05370 - 05374

  --0001010011111111    0001010100000000    0001010100000001    0001010100000010    0001010100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05375 - 05379

  --0001010100000100    0001010100000101    0001010100000110    0001010100000111    0001010100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05380 - 05384

  --0001010100001001    0001010100001010    0001010100001011    0001010100001100    0001010100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05385 - 05389

  --0001010100001110    0001010100001111    0001010100010000    0001010100010001    0001010100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05390 - 05394

  --0001010100010011    0001010100010100    0001010100010101    0001010100010110    0001010100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05395 - 05399

  --0001010100011000    0001010100011001    0001010100011010    0001010100011011    0001010100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05400 - 05404

  --0001010100011101    0001010100011110    0001010100011111    0001010100100000    0001010100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05405 - 05409

  --0001010100100010    0001010100100011    0001010100100100    0001010100100101    0001010100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05410 - 05414

  --0001010100100111    0001010100101000    0001010100101001    0001010100101010    0001010100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05415 - 05419

  --0001010100101100    0001010100101101    0001010100101110    0001010100101111    0001010100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05420 - 05424

  --0001010100110001    0001010100110010    0001010100110011    0001010100110100    0001010100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05425 - 05429

  --0001010100110110    0001010100110111    0001010100111000    0001010100111001    0001010100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05430 - 05434

  --0001010100111011    0001010100111100    0001010100111101    0001010100111110    0001010100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05435 - 05439

  --0001010101000000    0001010101000001    0001010101000010    0001010101000011    0001010101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05440 - 05444

  --0001010101000101    0001010101000110    0001010101000111    0001010101001000    0001010101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05445 - 05449

  --0001010101001010    0001010101001011    0001010101001100    0001010101001101    0001010101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05450 - 05454

  --0001010101001111    0001010101010000    0001010101010001    0001010101010010    0001010101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05455 - 05459

  --0001010101010100    0001010101010101    0001010101010110    0001010101010111    0001010101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05460 - 05464

  --0001010101011001    0001010101011010    0001010101011011    0001010101011100    0001010101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05465 - 05469

  --0001010101011110    0001010101011111    0001010101100000    0001010101100001    0001010101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05470 - 05474

  --0001010101100011    0001010101100100    0001010101100101    0001010101100110    0001010101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05475 - 05479

  --0001010101101000    0001010101101001    0001010101101010    0001010101101011    0001010101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05480 - 05484

  --0001010101101101    0001010101101110    0001010101101111    0001010101110000    0001010101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05485 - 05489

  --0001010101110010    0001010101110011    0001010101110100    0001010101110101    0001010101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05490 - 05494

  --0001010101110111    0001010101111000    0001010101111001    0001010101111010    0001010101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05495 - 05499

  --0001010101111100    0001010101111101    0001010101111110    0001010101111111    0001010110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05500 - 05504

  --0001010110000001    0001010110000010    0001010110000011    0001010110000100    0001010110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05505 - 05509

  --0001010110000110    0001010110000111    0001010110001000    0001010110001001    0001010110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05510 - 05514

  --0001010110001011    0001010110001100    0001010110001101    0001010110001110    0001010110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05515 - 05519

  --0001010110010000    0001010110010001    0001010110010010    0001010110010011    0001010110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05520 - 05524

  --0001010110010101    0001010110010110    0001010110010111    0001010110011000    0001010110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05525 - 05529

  --0001010110011010    0001010110011011    0001010110011100    0001010110011101    0001010110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05530 - 05534

  --0001010110011111    0001010110100000    0001010110100001    0001010110100010    0001010110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05535 - 05539

  --0001010110100100    0001010110100101    0001010110100110    0001010110100111    0001010110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05540 - 05544

  --0001010110101001    0001010110101010    0001010110101011    0001010110101100    0001010110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05545 - 05549

  --0001010110101110    0001010110101111    0001010110110000    0001010110110001    0001010110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05550 - 05554

  --0001010110110011    0001010110110100    0001010110110101    0001010110110110    0001010110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05555 - 05559

  --0001010110111000    0001010110111001    0001010110111010    0001010110111011    0001010110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05560 - 05564

  --0001010110111101    0001010110111110    0001010110111111    0001010111000000    0001010111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05565 - 05569

  --0001010111000010    0001010111000011    0001010111000100    0001010111000101    0001010111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05570 - 05574

  --0001010111000111    0001010111001000    0001010111001001    0001010111001010    0001010111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05575 - 05579

  --0001010111001100    0001010111001101    0001010111001110    0001010111001111    0001010111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05580 - 05584

  --0001010111010001    0001010111010010    0001010111010011    0001010111010100    0001010111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05585 - 05589

  --0001010111010110    0001010111010111    0001010111011000    0001010111011001    0001010111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05590 - 05594

  --0001010111011011    0001010111011100    0001010111011101    0001010111011110    0001010111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05595 - 05599

  --0001010111100000    0001010111100001    0001010111100010    0001010111100011    0001010111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05600 - 05604

  --0001010111100101    0001010111100110    0001010111100111    0001010111101000    0001010111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05605 - 05609

  --0001010111101010    0001010111101011    0001010111101100    0001010111101101    0001010111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05610 - 05614

  --0001010111101111    0001010111110000    0001010111110001    0001010111110010    0001010111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05615 - 05619

  --0001010111110100    0001010111110101    0001010111110110    0001010111110111    0001010111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05620 - 05624

  --0001010111111001    0001010111111010    0001010111111011    0001010111111100    0001010111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05625 - 05629

  --0001010111111110    0001010111111111    0001011000000000    0001011000000001    0001011000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05630 - 05634

  --0001011000000011    0001011000000100    0001011000000101    0001011000000110    0001011000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05635 - 05639

  --0001011000001000    0001011000001001    0001011000001010    0001011000001011    0001011000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05640 - 05644

  --0001011000001101    0001011000001110    0001011000001111    0001011000010000    0001011000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05645 - 05649

  --0001011000010010    0001011000010011    0001011000010100    0001011000010101    0001011000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05650 - 05654

  --0001011000010111    0001011000011000    0001011000011001    0001011000011010    0001011000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05655 - 05659

  --0001011000011100    0001011000011101    0001011000011110    0001011000011111    0001011000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05660 - 05664

  --0001011000100001    0001011000100010    0001011000100011    0001011000100100    0001011000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05665 - 05669

  --0001011000100110    0001011000100111    0001011000101000    0001011000101001    0001011000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05670 - 05674

  --0001011000101011    0001011000101100    0001011000101101    0001011000101110    0001011000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05675 - 05679

  --0001011000110000    0001011000110001    0001011000110010    0001011000110011    0001011000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05680 - 05684

  --0001011000110101    0001011000110110    0001011000110111    0001011000111000    0001011000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05685 - 05689

  --0001011000111010    0001011000111011    0001011000111100    0001011000111101    0001011000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05690 - 05694

  --0001011000111111    0001011001000000    0001011001000001    0001011001000010    0001011001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05695 - 05699

  --0001011001000100    0001011001000101    0001011001000110    0001011001000111    0001011001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05700 - 05704

  --0001011001001001    0001011001001010    0001011001001011    0001011001001100    0001011001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05705 - 05709

  --0001011001001110    0001011001001111    0001011001010000    0001011001010001    0001011001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05710 - 05714

  --0001011001010011    0001011001010100    0001011001010101    0001011001010110    0001011001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05715 - 05719

  --0001011001011000    0001011001011001    0001011001011010    0001011001011011    0001011001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05720 - 05724

  --0001011001011101    0001011001011110    0001011001011111    0001011001100000    0001011001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05725 - 05729

  --0001011001100010    0001011001100011    0001011001100100    0001011001100101    0001011001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05730 - 05734

  --0001011001100111    0001011001101000    0001011001101001    0001011001101010    0001011001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05735 - 05739

  --0001011001101100    0001011001101101    0001011001101110    0001011001101111    0001011001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05740 - 05744

  --0001011001110001    0001011001110010    0001011001110011    0001011001110100    0001011001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05745 - 05749

  --0001011001110110    0001011001110111    0001011001111000    0001011001111001    0001011001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05750 - 05754

  --0001011001111011    0001011001111100    0001011001111101    0001011001111110    0001011001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05755 - 05759

  --0001011010000000    0001011010000001    0001011010000010    0001011010000011    0001011010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05760 - 05764

  --0001011010000101    0001011010000110    0001011010000111    0001011010001000    0001011010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05765 - 05769

  --0001011010001010    0001011010001011    0001011010001100    0001011010001101    0001011010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05770 - 05774

  --0001011010001111    0001011010010000    0001011010010001    0001011010010010    0001011010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05775 - 05779

  --0001011010010100    0001011010010101    0001011010010110    0001011010010111    0001011010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05780 - 05784

  --0001011010011001    0001011010011010    0001011010011011    0001011010011100    0001011010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05785 - 05789

  --0001011010011110    0001011010011111    0001011010100000    0001011010100001    0001011010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05790 - 05794

  --0001011010100011    0001011010100100    0001011010100101    0001011010100110    0001011010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05795 - 05799

  --0001011010101000    0001011010101001    0001011010101010    0001011010101011    0001011010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05800 - 05804

  --0001011010101101    0001011010101110    0001011010101111    0001011010110000    0001011010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05805 - 05809

  --0001011010110010    0001011010110011    0001011010110100    0001011010110101    0001011010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05810 - 05814

  --0001011010110111    0001011010111000    0001011010111001    0001011010111010    0001011010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05815 - 05819

  --0001011010111100    0001011010111101    0001011010111110    0001011010111111    0001011011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05820 - 05824

  --0001011011000001    0001011011000010    0001011011000011    0001011011000100    0001011011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05825 - 05829

  --0001011011000110    0001011011000111    0001011011001000    0001011011001001    0001011011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05830 - 05834

  --0001011011001011    0001011011001100    0001011011001101    0001011011001110    0001011011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05835 - 05839

  --0001011011010000    0001011011010001    0001011011010010    0001011011010011    0001011011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05840 - 05844

  --0001011011010101    0001011011010110    0001011011010111    0001011011011000    0001011011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05845 - 05849

  --0001011011011010    0001011011011011    0001011011011100    0001011011011101    0001011011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05850 - 05854

  --0001011011011111    0001011011100000    0001011011100001    0001011011100010    0001011011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05855 - 05859

  --0001011011100100    0001011011100101    0001011011100110    0001011011100111    0001011011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05860 - 05864

  --0001011011101001    0001011011101010    0001011011101011    0001011011101100    0001011011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05865 - 05869

  --0001011011101110    0001011011101111    0001011011110000    0001011011110001    0001011011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05870 - 05874

  --0001011011110011    0001011011110100    0001011011110101    0001011011110110    0001011011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05875 - 05879

  --0001011011111000    0001011011111001    0001011011111010    0001011011111011    0001011011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05880 - 05884

  --0001011011111101    0001011011111110    0001011011111111    0001011100000000    0001011100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05885 - 05889

  --0001011100000010    0001011100000011    0001011100000100    0001011100000101    0001011100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05890 - 05894

  --0001011100000111    0001011100001000    0001011100001001    0001011100001010    0001011100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05895 - 05899

  --0001011100001100    0001011100001101    0001011100001110    0001011100001111    0001011100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05900 - 05904

  --0001011100010001    0001011100010010    0001011100010011    0001011100010100    0001011100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05905 - 05909

  --0001011100010110    0001011100010111    0001011100011000    0001011100011001    0001011100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05910 - 05914

  --0001011100011011    0001011100011100    0001011100011101    0001011100011110    0001011100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05915 - 05919

  --0001011100100000    0001011100100001    0001011100100010    0001011100100011    0001011100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05920 - 05924

  --0001011100100101    0001011100100110    0001011100100111    0001011100101000    0001011100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05925 - 05929

  --0001011100101010    0001011100101011    0001011100101100    0001011100101101    0001011100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05930 - 05934

  --0001011100101111    0001011100110000    0001011100110001    0001011100110010    0001011100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05935 - 05939

  --0001011100110100    0001011100110101    0001011100110110    0001011100110111    0001011100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05940 - 05944

  --0001011100111001    0001011100111010    0001011100111011    0001011100111100    0001011100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05945 - 05949

  --0001011100111110    0001011100111111    0001011101000000    0001011101000001    0001011101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05950 - 05954

  --0001011101000011    0001011101000100    0001011101000101    0001011101000110    0001011101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05955 - 05959

  --0001011101001000    0001011101001001    0001011101001010    0001011101001011    0001011101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05960 - 05964

  --0001011101001101    0001011101001110    0001011101001111    0001011101010000    0001011101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05965 - 05969

  --0001011101010010    0001011101010011    0001011101010100    0001011101010101    0001011101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05970 - 05974

  --0001011101010111    0001011101011000    0001011101011001    0001011101011010    0001011101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05975 - 05979

  --0001011101011100    0001011101011101    0001011101011110    0001011101011111    0001011101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05980 - 05984

  --0001011101100001    0001011101100010    0001011101100011    0001011101100100    0001011101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05985 - 05989

  --0001011101100110    0001011101100111    0001011101101000    0001011101101001    0001011101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05990 - 05994

  --0001011101101011    0001011101101100    0001011101101101    0001011101101110    0001011101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 05995 - 05999

  --0001011101110000    0001011101110001    0001011101110010    0001011101110011    0001011101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06000 - 06004

  --0001011101110101    0001011101110110    0001011101110111    0001011101111000    0001011101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06005 - 06009

  --0001011101111010    0001011101111011    0001011101111100    0001011101111101    0001011101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06010 - 06014

  --0001011101111111    0001011110000000    0001011110000001    0001011110000010    0001011110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06015 - 06019

  --0001011110000100    0001011110000101    0001011110000110    0001011110000111    0001011110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06020 - 06024

  --0001011110001001    0001011110001010    0001011110001011    0001011110001100    0001011110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06025 - 06029

  --0001011110001110    0001011110001111    0001011110010000    0001011110010001    0001011110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06030 - 06034

  --0001011110010011    0001011110010100    0001011110010101    0001011110010110    0001011110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06035 - 06039

  --0001011110011000    0001011110011001    0001011110011010    0001011110011011    0001011110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06040 - 06044

  --0001011110011101    0001011110011110    0001011110011111    0001011110100000    0001011110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06045 - 06049

  --0001011110100010    0001011110100011    0001011110100100    0001011110100101    0001011110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06050 - 06054

  --0001011110100111    0001011110101000    0001011110101001    0001011110101010    0001011110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06055 - 06059

  --0001011110101100    0001011110101101    0001011110101110    0001011110101111    0001011110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06060 - 06064

  --0001011110110001    0001011110110010    0001011110110011    0001011110110100    0001011110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06065 - 06069

  --0001011110110110    0001011110110111    0001011110111000    0001011110111001    0001011110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06070 - 06074

  --0001011110111011    0001011110111100    0001011110111101    0001011110111110    0001011110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06075 - 06079

  --0001011111000000    0001011111000001    0001011111000010    0001011111000011    0001011111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06080 - 06084

  --0001011111000101    0001011111000110    0001011111000111    0001011111001000    0001011111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06085 - 06089

  --0001011111001010    0001011111001011    0001011111001100    0001011111001101    0001011111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06090 - 06094

  --0001011111001111    0001011111010000    0001011111010001    0001011111010010    0001011111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06095 - 06099

  --0001011111010100    0001011111010101    0001011111010110    0001011111010111    0001011111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06100 - 06104

  --0001011111011001    0001011111011010    0001011111011011    0001011111011100    0001011111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06105 - 06109

  --0001011111011110    0001011111011111    0001011111100000    0001011111100001    0001011111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06110 - 06114

  --0001011111100011    0001011111100100    0001011111100101    0001011111100110    0001011111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06115 - 06119

  --0001011111101000    0001011111101001    0001011111101010    0001011111101011    0001011111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06120 - 06124

  --0001011111101101    0001011111101110    0001011111101111    0001011111110000    0001011111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06125 - 06129

  --0001011111110010    0001011111110011    0001011111110100    0001011111110101    0001011111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06130 - 06134

  --0001011111110111    0001011111111000    0001011111111001    0001011111111010    0001011111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06135 - 06139

  --0001011111111100    0001011111111101    0001011111111110    0001011111111111    0001100000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06140 - 06144

  --0001100000000001    0001100000000010    0001100000000011    0001100000000100    0001100000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06145 - 06149

  --0001100000000110    0001100000000111    0001100000001000    0001100000001001    0001100000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06150 - 06154

  --0001100000001011    0001100000001100    0001100000001101    0001100000001110    0001100000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06155 - 06159

  --0001100000010000    0001100000010001    0001100000010010    0001100000010011    0001100000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06160 - 06164

  --0001100000010101    0001100000010110    0001100000010111    0001100000011000    0001100000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06165 - 06169

  --0001100000011010    0001100000011011    0001100000011100    0001100000011101    0001100000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06170 - 06174

  --0001100000011111    0001100000100000    0001100000100001    0001100000100010    0001100000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06175 - 06179

  --0001100000100100    0001100000100101    0001100000100110    0001100000100111    0001100000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06180 - 06184

  --0001100000101001    0001100000101010    0001100000101011    0001100000101100    0001100000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06185 - 06189

  --0001100000101110    0001100000101111    0001100000110000    0001100000110001    0001100000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06190 - 06194

  --0001100000110011    0001100000110100    0001100000110101    0001100000110110    0001100000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06195 - 06199

  --0001100000111000    0001100000111001    0001100000111010    0001100000111011    0001100000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06200 - 06204

  --0001100000111101    0001100000111110    0001100000111111    0001100001000000    0001100001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06205 - 06209

  --0001100001000010    0001100001000011    0001100001000100    0001100001000101    0001100001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06210 - 06214

  --0001100001000111    0001100001001000    0001100001001001    0001100001001010    0001100001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06215 - 06219

  --0001100001001100    0001100001001101    0001100001001110    0001100001001111    0001100001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06220 - 06224

  --0001100001010001    0001100001010010    0001100001010011    0001100001010100    0001100001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06225 - 06229

  --0001100001010110    0001100001010111    0001100001011000    0001100001011001    0001100001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06230 - 06234

  --0001100001011011    0001100001011100    0001100001011101    0001100001011110    0001100001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06235 - 06239

  --0001100001100000    0001100001100001    0001100001100010    0001100001100011    0001100001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06240 - 06244

  --0001100001100101    0001100001100110    0001100001100111    0001100001101000    0001100001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06245 - 06249

  --0001100001101010    0001100001101011    0001100001101100    0001100001101101    0001100001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06250 - 06254

  --0001100001101111    0001100001110000    0001100001110001    0001100001110010    0001100001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06255 - 06259

  --0001100001110100    0001100001110101    0001100001110110    0001100001110111    0001100001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06260 - 06264

  --0001100001111001    0001100001111010    0001100001111011    0001100001111100    0001100001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06265 - 06269

  --0001100001111110    0001100001111111    0001100010000000    0001100010000001    0001100010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06270 - 06274

  --0001100010000011    0001100010000100    0001100010000101    0001100010000110    0001100010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06275 - 06279

  --0001100010001000    0001100010001001    0001100010001010    0001100010001011    0001100010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06280 - 06284

  --0001100010001101    0001100010001110    0001100010001111    0001100010010000    0001100010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06285 - 06289

  --0001100010010010    0001100010010011    0001100010010100    0001100010010101    0001100010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06290 - 06294

  --0001100010010111    0001100010011000    0001100010011001    0001100010011010    0001100010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06295 - 06299

  --0001100010011100    0001100010011101    0001100010011110    0001100010011111    0001100010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06300 - 06304

  --0001100010100001    0001100010100010    0001100010100011    0001100010100100    0001100010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06305 - 06309

  --0001100010100110    0001100010100111    0001100010101000    0001100010101001    0001100010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06310 - 06314

  --0001100010101011    0001100010101100    0001100010101101    0001100010101110    0001100010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06315 - 06319

  --0001100010110000    0001100010110001    0001100010110010    0001100010110011    0001100010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06320 - 06324

  --0001100010110101    0001100010110110    0001100010110111    0001100010111000    0001100010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06325 - 06329

  --0001100010111010    0001100010111011    0001100010111100    0001100010111101    0001100010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06330 - 06334

  --0001100010111111    0001100011000000    0001100011000001    0001100011000010    0001100011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06335 - 06339

  --0001100011000100    0001100011000101    0001100011000110    0001100011000111    0001100011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06340 - 06344

  --0001100011001001    0001100011001010    0001100011001011    0001100011001100    0001100011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06345 - 06349

  --0001100011001110    0001100011001111    0001100011010000    0001100011010001    0001100011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06350 - 06354

  --0001100011010011    0001100011010100    0001100011010101    0001100011010110    0001100011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06355 - 06359

  --0001100011011000    0001100011011001    0001100011011010    0001100011011011    0001100011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06360 - 06364

  --0001100011011101    0001100011011110    0001100011011111    0001100011100000    0001100011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06365 - 06369

  --0001100011100010    0001100011100011    0001100011100100    0001100011100101    0001100011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06370 - 06374

  --0001100011100111    0001100011101000    0001100011101001    0001100011101010    0001100011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06375 - 06379

  --0001100011101100    0001100011101101    0001100011101110    0001100011101111    0001100011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06380 - 06384

  --0001100011110001    0001100011110010    0001100011110011    0001100011110100    0001100011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06385 - 06389

  --0001100011110110    0001100011110111    0001100011111000    0001100011111001    0001100011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06390 - 06394

  --0001100011111011    0001100011111100    0001100011111101    0001100011111110    0001100011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06395 - 06399

  --0001100100000000    0001100100000001    0001100100000010    0001100100000011    0001100100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06400 - 06404

  --0001100100000101    0001100100000110    0001100100000111    0001100100001000    0001100100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06405 - 06409

  --0001100100001010    0001100100001011    0001100100001100    0001100100001101    0001100100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06410 - 06414

  --0001100100001111    0001100100010000    0001100100010001    0001100100010010    0001100100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06415 - 06419

  --0001100100010100    0001100100010101    0001100100010110    0001100100010111    0001100100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06420 - 06424

  --0001100100011001    0001100100011010    0001100100011011    0001100100011100    0001100100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06425 - 06429

  --0001100100011110    0001100100011111    0001100100100000    0001100100100001    0001100100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06430 - 06434

  --0001100100100011    0001100100100100    0001100100100101    0001100100100110    0001100100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06435 - 06439

  --0001100100101000    0001100100101001    0001100100101010    0001100100101011    0001100100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06440 - 06444

  --0001100100101101    0001100100101110    0001100100101111    0001100100110000    0001100100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06445 - 06449

  --0001100100110010    0001100100110011    0001100100110100    0001100100110101    0001100100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06450 - 06454

  --0001100100110111    0001100100111000    0001100100111001    0001100100111010    0001100100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06455 - 06459

  --0001100100111100    0001100100111101    0001100100111110    0001100100111111    0001100101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06460 - 06464

  --0001100101000001    0001100101000010    0001100101000011    0001100101000100    0001100101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06465 - 06469

  --0001100101000110    0001100101000111    0001100101001000    0001100101001001    0001100101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06470 - 06474

  --0001100101001011    0001100101001100    0001100101001101    0001100101001110    0001100101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06475 - 06479

  --0001100101010000    0001100101010001    0001100101010010    0001100101010011    0001100101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06480 - 06484

  --0001100101010101    0001100101010110    0001100101010111    0001100101011000    0001100101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06485 - 06489

  --0001100101011010    0001100101011011    0001100101011100    0001100101011101    0001100101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06490 - 06494

  --0001100101011111    0001100101100000    0001100101100001    0001100101100010    0001100101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06495 - 06499

  --0001100101100100    0001100101100101    0001100101100110    0001100101100111    0001100101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06500 - 06504

  --0001100101101001    0001100101101010    0001100101101011    0001100101101100    0001100101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06505 - 06509

  --0001100101101110    0001100101101111    0001100101110000    0001100101110001    0001100101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06510 - 06514

  --0001100101110011    0001100101110100    0001100101110101    0001100101110110    0001100101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06515 - 06519

  --0001100101111000    0001100101111001    0001100101111010    0001100101111011    0001100101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06520 - 06524

  --0001100101111101    0001100101111110    0001100101111111    0001100110000000    0001100110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06525 - 06529

  --0001100110000010    0001100110000011    0001100110000100    0001100110000101    0001100110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06530 - 06534

  --0001100110000111    0001100110001000    0001100110001001    0001100110001010    0001100110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06535 - 06539

  --0001100110001100    0001100110001101    0001100110001110    0001100110001111    0001100110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06540 - 06544

  --0001100110010001    0001100110010010    0001100110010011    0001100110010100    0001100110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06545 - 06549

  --0001100110010110    0001100110010111    0001100110011000    0001100110011001    0001100110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06550 - 06554

  --0001100110011011    0001100110011100    0001100110011101    0001100110011110    0001100110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06555 - 06559

  --0001100110100000    0001100110100001    0001100110100010    0001100110100011    0001100110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06560 - 06564

  --0001100110100101    0001100110100110    0001100110100111    0001100110101000    0001100110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06565 - 06569

  --0001100110101010    0001100110101011    0001100110101100    0001100110101101    0001100110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06570 - 06574

  --0001100110101111    0001100110110000    0001100110110001    0001100110110010    0001100110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06575 - 06579

  --0001100110110100    0001100110110101    0001100110110110    0001100110110111    0001100110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06580 - 06584

  --0001100110111001    0001100110111010    0001100110111011    0001100110111100    0001100110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06585 - 06589

  --0001100110111110    0001100110111111    0001100111000000    0001100111000001    0001100111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06590 - 06594

  --0001100111000011    0001100111000100    0001100111000101    0001100111000110    0001100111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06595 - 06599

  --0001100111001000    0001100111001001    0001100111001010    0001100111001011    0001100111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06600 - 06604

  --0001100111001101    0001100111001110    0001100111001111    0001100111010000    0001100111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06605 - 06609

  --0001100111010010    0001100111010011    0001100111010100    0001100111010101    0001100111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06610 - 06614

  --0001100111010111    0001100111011000    0001100111011001    0001100111011010    0001100111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06615 - 06619

  --0001100111011100    0001100111011101    0001100111011110    0001100111011111    0001100111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06620 - 06624

  --0001100111100001    0001100111100010    0001100111100011    0001100111100100    0001100111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06625 - 06629

  --0001100111100110    0001100111100111    0001100111101000    0001100111101001    0001100111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06630 - 06634

  --0001100111101011    0001100111101100    0001100111101101    0001100111101110    0001100111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06635 - 06639

  --0001100111110000    0001100111110001    0001100111110010    0001100111110011    0001100111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06640 - 06644

  --0001100111110101    0001100111110110    0001100111110111    0001100111111000    0001100111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06645 - 06649

  --0001100111111010    0001100111111011    0001100111111100    0001100111111101    0001100111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06650 - 06654

  --0001100111111111    0001101000000000    0001101000000001    0001101000000010    0001101000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06655 - 06659

  --0001101000000100    0001101000000101    0001101000000110    0001101000000111    0001101000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06660 - 06664

  --0001101000001001    0001101000001010    0001101000001011    0001101000001100    0001101000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06665 - 06669

  --0001101000001110    0001101000001111    0001101000010000    0001101000010001    0001101000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06670 - 06674

  --0001101000010011    0001101000010100    0001101000010101    0001101000010110    0001101000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06675 - 06679

  --0001101000011000    0001101000011001    0001101000011010    0001101000011011    0001101000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06680 - 06684

  --0001101000011101    0001101000011110    0001101000011111    0001101000100000    0001101000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06685 - 06689

  --0001101000100010    0001101000100011    0001101000100100    0001101000100101    0001101000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06690 - 06694

  --0001101000100111    0001101000101000    0001101000101001    0001101000101010    0001101000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06695 - 06699

  --0001101000101100    0001101000101101    0001101000101110    0001101000101111    0001101000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06700 - 06704

  --0001101000110001    0001101000110010    0001101000110011    0001101000110100    0001101000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06705 - 06709

  --0001101000110110    0001101000110111    0001101000111000    0001101000111001    0001101000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06710 - 06714

  --0001101000111011    0001101000111100    0001101000111101    0001101000111110    0001101000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06715 - 06719

  --0001101001000000    0001101001000001    0001101001000010    0001101001000011    0001101001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06720 - 06724

  --0001101001000101    0001101001000110    0001101001000111    0001101001001000    0001101001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06725 - 06729

  --0001101001001010    0001101001001011    0001101001001100    0001101001001101    0001101001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06730 - 06734

  --0001101001001111    0001101001010000    0001101001010001    0001101001010010    0001101001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06735 - 06739

  --0001101001010100    0001101001010101    0001101001010110    0001101001010111    0001101001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06740 - 06744

  --0001101001011001    0001101001011010    0001101001011011    0001101001011100    0001101001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06745 - 06749

  --0001101001011110    0001101001011111    0001101001100000    0001101001100001    0001101001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06750 - 06754

  --0001101001100011    0001101001100100    0001101001100101    0001101001100110    0001101001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06755 - 06759

  --0001101001101000    0001101001101001    0001101001101010    0001101001101011    0001101001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06760 - 06764

  --0001101001101101    0001101001101110    0001101001101111    0001101001110000    0001101001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06765 - 06769

  --0001101001110010    0001101001110011    0001101001110100    0001101001110101    0001101001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06770 - 06774

  --0001101001110111    0001101001111000    0001101001111001    0001101001111010    0001101001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06775 - 06779

  --0001101001111100    0001101001111101    0001101001111110    0001101001111111    0001101010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06780 - 06784

  --0001101010000001    0001101010000010    0001101010000011    0001101010000100    0001101010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06785 - 06789

  --0001101010000110    0001101010000111    0001101010001000    0001101010001001    0001101010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06790 - 06794

  --0001101010001011    0001101010001100    0001101010001101    0001101010001110    0001101010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06795 - 06799

  --0001101010010000    0001101010010001    0001101010010010    0001101010010011    0001101010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06800 - 06804

  --0001101010010101    0001101010010110    0001101010010111    0001101010011000    0001101010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06805 - 06809

  --0001101010011010    0001101010011011    0001101010011100    0001101010011101    0001101010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06810 - 06814

  --0001101010011111    0001101010100000    0001101010100001    0001101010100010    0001101010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06815 - 06819

  --0001101010100100    0001101010100101    0001101010100110    0001101010100111    0001101010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06820 - 06824

  --0001101010101001    0001101010101010    0001101010101011    0001101010101100    0001101010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06825 - 06829

  --0001101010101110    0001101010101111    0001101010110000    0001101010110001    0001101010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06830 - 06834

  --0001101010110011    0001101010110100    0001101010110101    0001101010110110    0001101010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06835 - 06839

  --0001101010111000    0001101010111001    0001101010111010    0001101010111011    0001101010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06840 - 06844

  --0001101010111101    0001101010111110    0001101010111111    0001101011000000    0001101011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06845 - 06849

  --0001101011000010    0001101011000011    0001101011000100    0001101011000101    0001101011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06850 - 06854

  --0001101011000111    0001101011001000    0001101011001001    0001101011001010    0001101011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06855 - 06859

  --0001101011001100    0001101011001101    0001101011001110    0001101011001111    0001101011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06860 - 06864

  --0001101011010001    0001101011010010    0001101011010011    0001101011010100    0001101011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06865 - 06869

  --0001101011010110    0001101011010111    0001101011011000    0001101011011001    0001101011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06870 - 06874

  --0001101011011011    0001101011011100    0001101011011101    0001101011011110    0001101011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06875 - 06879

  --0001101011100000    0001101011100001    0001101011100010    0001101011100011    0001101011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06880 - 06884

  --0001101011100101    0001101011100110    0001101011100111    0001101011101000    0001101011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06885 - 06889

  --0001101011101010    0001101011101011    0001101011101100    0001101011101101    0001101011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06890 - 06894

  --0001101011101111    0001101011110000    0001101011110001    0001101011110010    0001101011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06895 - 06899

  --0001101011110100    0001101011110101    0001101011110110    0001101011110111    0001101011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06900 - 06904

  --0001101011111001    0001101011111010    0001101011111011    0001101011111100    0001101011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06905 - 06909

  --0001101011111110    0001101011111111    0001101100000000    0001101100000001    0001101100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06910 - 06914

  --0001101100000011    0001101100000100    0001101100000101    0001101100000110    0001101100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06915 - 06919

  --0001101100001000    0001101100001001    0001101100001010    0001101100001011    0001101100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06920 - 06924

  --0001101100001101    0001101100001110    0001101100001111    0001101100010000    0001101100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06925 - 06929

  --0001101100010010    0001101100010011    0001101100010100    0001101100010101    0001101100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06930 - 06934

  --0001101100010111    0001101100011000    0001101100011001    0001101100011010    0001101100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06935 - 06939

  --0001101100011100    0001101100011101    0001101100011110    0001101100011111    0001101100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06940 - 06944

  --0001101100100001    0001101100100010    0001101100100011    0001101100100100    0001101100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06945 - 06949

  --0001101100100110    0001101100100111    0001101100101000    0001101100101001    0001101100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06950 - 06954

  --0001101100101011    0001101100101100    0001101100101101    0001101100101110    0001101100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06955 - 06959

  --0001101100110000    0001101100110001    0001101100110010    0001101100110011    0001101100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06960 - 06964

  --0001101100110101    0001101100110110    0001101100110111    0001101100111000    0001101100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06965 - 06969

  --0001101100111010    0001101100111011    0001101100111100    0001101100111101    0001101100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06970 - 06974

  --0001101100111111    0001101101000000    0001101101000001    0001101101000010    0001101101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06975 - 06979

  --0001101101000100    0001101101000101    0001101101000110    0001101101000111    0001101101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06980 - 06984

  --0001101101001001    0001101101001010    0001101101001011    0001101101001100    0001101101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06985 - 06989

  --0001101101001110    0001101101001111    0001101101010000    0001101101010001    0001101101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06990 - 06994

  --0001101101010011    0001101101010100    0001101101010101    0001101101010110    0001101101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 06995 - 06999

  --0001101101011000    0001101101011001    0001101101011010    0001101101011011    0001101101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07000 - 07004

  --0001101101011101    0001101101011110    0001101101011111    0001101101100000    0001101101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07005 - 07009

  --0001101101100010    0001101101100011    0001101101100100    0001101101100101    0001101101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07010 - 07014

  --0001101101100111    0001101101101000    0001101101101001    0001101101101010    0001101101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07015 - 07019

  --0001101101101100    0001101101101101    0001101101101110    0001101101101111    0001101101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07020 - 07024

  --0001101101110001    0001101101110010    0001101101110011    0001101101110100    0001101101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07025 - 07029

  --0001101101110110    0001101101110111    0001101101111000    0001101101111001    0001101101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07030 - 07034

  --0001101101111011    0001101101111100    0001101101111101    0001101101111110    0001101101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07035 - 07039

  --0001101110000000    0001101110000001    0001101110000010    0001101110000011    0001101110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07040 - 07044

  --0001101110000101    0001101110000110    0001101110000111    0001101110001000    0001101110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07045 - 07049

  --0001101110001010    0001101110001011    0001101110001100    0001101110001101    0001101110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07050 - 07054

  --0001101110001111    0001101110010000    0001101110010001    0001101110010010    0001101110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07055 - 07059

  --0001101110010100    0001101110010101    0001101110010110    0001101110010111    0001101110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07060 - 07064

  --0001101110011001    0001101110011010    0001101110011011    0001101110011100    0001101110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07065 - 07069

  --0001101110011110    0001101110011111    0001101110100000    0001101110100001    0001101110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07070 - 07074

  --0001101110100011    0001101110100100    0001101110100101    0001101110100110    0001101110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07075 - 07079

  --0001101110101000    0001101110101001    0001101110101010    0001101110101011    0001101110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07080 - 07084

  --0001101110101101    0001101110101110    0001101110101111    0001101110110000    0001101110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07085 - 07089

  --0001101110110010    0001101110110011    0001101110110100    0001101110110101    0001101110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07090 - 07094

  --0001101110110111    0001101110111000    0001101110111001    0001101110111010    0001101110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07095 - 07099

  --0001101110111100    0001101110111101    0001101110111110    0001101110111111    0001101111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07100 - 07104

  --0001101111000001    0001101111000010    0001101111000011    0001101111000100    0001101111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07105 - 07109

  --0001101111000110    0001101111000111    0001101111001000    0001101111001001    0001101111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07110 - 07114

  --0001101111001011    0001101111001100    0001101111001101    0001101111001110    0001101111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07115 - 07119

  --0001101111010000    0001101111010001    0001101111010010    0001101111010011    0001101111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07120 - 07124

  --0001101111010101    0001101111010110    0001101111010111    0001101111011000    0001101111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07125 - 07129

  --0001101111011010    0001101111011011    0001101111011100    0001101111011101    0001101111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07130 - 07134

  --0001101111011111    0001101111100000    0001101111100001    0001101111100010    0001101111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07135 - 07139

  --0001101111100100    0001101111100101    0001101111100110    0001101111100111    0001101111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07140 - 07144

  --0001101111101001    0001101111101010    0001101111101011    0001101111101100    0001101111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07145 - 07149

  --0001101111101110    0001101111101111    0001101111110000    0001101111110001    0001101111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07150 - 07154

  --0001101111110011    0001101111110100    0001101111110101    0001101111110110    0001101111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07155 - 07159

  --0001101111111000    0001101111111001    0001101111111010    0001101111111011    0001101111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07160 - 07164

  --0001101111111101    0001101111111110    0001101111111111    0001110000000000    0001110000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07165 - 07169

  --0001110000000010    0001110000000011    0001110000000100    0001110000000101    0001110000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07170 - 07174

  --0001110000000111    0001110000001000    0001110000001001    0001110000001010    0001110000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07175 - 07179

  --0001110000001100    0001110000001101    0001110000001110    0001110000001111    0001110000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07180 - 07184

  --0001110000010001    0001110000010010    0001110000010011    0001110000010100    0001110000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07185 - 07189

  --0001110000010110    0001110000010111    0001110000011000    0001110000011001    0001110000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07190 - 07194

  --0001110000011011    0001110000011100    0001110000011101    0001110000011110    0001110000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07195 - 07199

  --0001110000100000    0001110000100001    0001110000100010    0001110000100011    0001110000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07200 - 07204

  --0001110000100101    0001110000100110    0001110000100111    0001110000101000    0001110000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07205 - 07209

  --0001110000101010    0001110000101011    0001110000101100    0001110000101101    0001110000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07210 - 07214

  --0001110000101111    0001110000110000    0001110000110001    0001110000110010    0001110000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07215 - 07219

  --0001110000110100    0001110000110101    0001110000110110    0001110000110111    0001110000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07220 - 07224

  --0001110000111001    0001110000111010    0001110000111011    0001110000111100    0001110000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07225 - 07229

  --0001110000111110    0001110000111111    0001110001000000    0001110001000001    0001110001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07230 - 07234

  --0001110001000011    0001110001000100    0001110001000101    0001110001000110    0001110001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07235 - 07239

  --0001110001001000    0001110001001001    0001110001001010    0001110001001011    0001110001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07240 - 07244

  --0001110001001101    0001110001001110    0001110001001111    0001110001010000    0001110001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07245 - 07249

  --0001110001010010    0001110001010011    0001110001010100    0001110001010101    0001110001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07250 - 07254

  --0001110001010111    0001110001011000    0001110001011001    0001110001011010    0001110001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07255 - 07259

  --0001110001011100    0001110001011101    0001110001011110    0001110001011111    0001110001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07260 - 07264

  --0001110001100001    0001110001100010    0001110001100011    0001110001100100    0001110001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07265 - 07269

  --0001110001100110    0001110001100111    0001110001101000    0001110001101001    0001110001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07270 - 07274

  --0001110001101011    0001110001101100    0001110001101101    0001110001101110    0001110001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07275 - 07279

  --0001110001110000    0001110001110001    0001110001110010    0001110001110011    0001110001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07280 - 07284

  --0001110001110101    0001110001110110    0001110001110111    0001110001111000    0001110001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07285 - 07289

  --0001110001111010    0001110001111011    0001110001111100    0001110001111101    0001110001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07290 - 07294

  --0001110001111111    0001110010000000    0001110010000001    0001110010000010    0001110010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07295 - 07299

  --0001110010000100    0001110010000101    0001110010000110    0001110010000111    0001110010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07300 - 07304

  --0001110010001001    0001110010001010    0001110010001011    0001110010001100    0001110010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07305 - 07309

  --0001110010001110    0001110010001111    0001110010010000    0001110010010001    0001110010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07310 - 07314

  --0001110010010011    0001110010010100    0001110010010101    0001110010010110    0001110010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07315 - 07319

  --0001110010011000    0001110010011001    0001110010011010    0001110010011011    0001110010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07320 - 07324

  --0001110010011101    0001110010011110    0001110010011111    0001110010100000    0001110010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07325 - 07329

  --0001110010100010    0001110010100011    0001110010100100    0001110010100101    0001110010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07330 - 07334

  --0001110010100111    0001110010101000    0001110010101001    0001110010101010    0001110010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07335 - 07339

  --0001110010101100    0001110010101101    0001110010101110    0001110010101111    0001110010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07340 - 07344

  --0001110010110001    0001110010110010    0001110010110011    0001110010110100    0001110010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07345 - 07349

  --0001110010110110    0001110010110111    0001110010111000    0001110010111001    0001110010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07350 - 07354

  --0001110010111011    0001110010111100    0001110010111101    0001110010111110    0001110010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07355 - 07359

  --0001110011000000    0001110011000001    0001110011000010    0001110011000011    0001110011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07360 - 07364

  --0001110011000101    0001110011000110    0001110011000111    0001110011001000    0001110011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07365 - 07369

  --0001110011001010    0001110011001011    0001110011001100    0001110011001101    0001110011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07370 - 07374

  --0001110011001111    0001110011010000    0001110011010001    0001110011010010    0001110011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07375 - 07379

  --0001110011010100    0001110011010101    0001110011010110    0001110011010111    0001110011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07380 - 07384

  --0001110011011001    0001110011011010    0001110011011011    0001110011011100    0001110011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07385 - 07389

  --0001110011011110    0001110011011111    0001110011100000    0001110011100001    0001110011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07390 - 07394

  --0001110011100011    0001110011100100    0001110011100101    0001110011100110    0001110011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07395 - 07399

  --0001110011101000    0001110011101001    0001110011101010    0001110011101011    0001110011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07400 - 07404

  --0001110011101101    0001110011101110    0001110011101111    0001110011110000    0001110011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07405 - 07409

  --0001110011110010    0001110011110011    0001110011110100    0001110011110101    0001110011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07410 - 07414

  --0001110011110111    0001110011111000    0001110011111001    0001110011111010    0001110011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07415 - 07419

  --0001110011111100    0001110011111101    0001110011111110    0001110011111111    0001110100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07420 - 07424

  --0001110100000001    0001110100000010    0001110100000011    0001110100000100    0001110100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07425 - 07429

  --0001110100000110    0001110100000111    0001110100001000    0001110100001001    0001110100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07430 - 07434

  --0001110100001011    0001110100001100    0001110100001101    0001110100001110    0001110100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07435 - 07439

  --0001110100010000    0001110100010001    0001110100010010    0001110100010011    0001110100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07440 - 07444

  --0001110100010101    0001110100010110    0001110100010111    0001110100011000    0001110100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07445 - 07449

  --0001110100011010    0001110100011011    0001110100011100    0001110100011101    0001110100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07450 - 07454

  --0001110100011111    0001110100100000    0001110100100001    0001110100100010    0001110100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07455 - 07459

  --0001110100100100    0001110100100101    0001110100100110    0001110100100111    0001110100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07460 - 07464

  --0001110100101001    0001110100101010    0001110100101011    0001110100101100    0001110100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07465 - 07469

  --0001110100101110    0001110100101111    0001110100110000    0001110100110001    0001110100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07470 - 07474

  --0001110100110011    0001110100110100    0001110100110101    0001110100110110    0001110100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07475 - 07479

  --0001110100111000    0001110100111001    0001110100111010    0001110100111011    0001110100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07480 - 07484

  --0001110100111101    0001110100111110    0001110100111111    0001110101000000    0001110101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07485 - 07489

  --0001110101000010    0001110101000011    0001110101000100    0001110101000101    0001110101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07490 - 07494

  --0001110101000111    0001110101001000    0001110101001001    0001110101001010    0001110101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07495 - 07499

  --0001110101001100    0001110101001101    0001110101001110    0001110101001111    0001110101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07500 - 07504

  --0001110101010001    0001110101010010    0001110101010011    0001110101010100    0001110101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07505 - 07509

  --0001110101010110    0001110101010111    0001110101011000    0001110101011001    0001110101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07510 - 07514

  --0001110101011011    0001110101011100    0001110101011101    0001110101011110    0001110101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07515 - 07519

  --0001110101100000    0001110101100001    0001110101100010    0001110101100011    0001110101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07520 - 07524

  --0001110101100101    0001110101100110    0001110101100111    0001110101101000    0001110101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07525 - 07529

  --0001110101101010    0001110101101011    0001110101101100    0001110101101101    0001110101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07530 - 07534

  --0001110101101111    0001110101110000    0001110101110001    0001110101110010    0001110101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07535 - 07539

  --0001110101110100    0001110101110101    0001110101110110    0001110101110111    0001110101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07540 - 07544

  --0001110101111001    0001110101111010    0001110101111011    0001110101111100    0001110101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07545 - 07549

  --0001110101111110    0001110101111111    0001110110000000    0001110110000001    0001110110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07550 - 07554

  --0001110110000011    0001110110000100    0001110110000101    0001110110000110    0001110110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07555 - 07559

  --0001110110001000    0001110110001001    0001110110001010    0001110110001011    0001110110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07560 - 07564

  --0001110110001101    0001110110001110    0001110110001111    0001110110010000    0001110110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07565 - 07569

  --0001110110010010    0001110110010011    0001110110010100    0001110110010101    0001110110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07570 - 07574

  --0001110110010111    0001110110011000    0001110110011001    0001110110011010    0001110110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07575 - 07579

  --0001110110011100    0001110110011101    0001110110011110    0001110110011111    0001110110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07580 - 07584

  --0001110110100001    0001110110100010    0001110110100011    0001110110100100    0001110110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07585 - 07589

  --0001110110100110    0001110110100111    0001110110101000    0001110110101001    0001110110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07590 - 07594

  --0001110110101011    0001110110101100    0001110110101101    0001110110101110    0001110110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07595 - 07599

  --0001110110110000    0001110110110001    0001110110110010    0001110110110011    0001110110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07600 - 07604

  --0001110110110101    0001110110110110    0001110110110111    0001110110111000    0001110110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07605 - 07609

  --0001110110111010    0001110110111011    0001110110111100    0001110110111101    0001110110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07610 - 07614

  --0001110110111111    0001110111000000    0001110111000001    0001110111000010    0001110111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07615 - 07619

  --0001110111000100    0001110111000101    0001110111000110    0001110111000111    0001110111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07620 - 07624

  --0001110111001001    0001110111001010    0001110111001011    0001110111001100    0001110111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07625 - 07629

  --0001110111001110    0001110111001111    0001110111010000    0001110111010001    0001110111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07630 - 07634

  --0001110111010011    0001110111010100    0001110111010101    0001110111010110    0001110111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07635 - 07639

  --0001110111011000    0001110111011001    0001110111011010    0001110111011011    0001110111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07640 - 07644

  --0001110111011101    0001110111011110    0001110111011111    0001110111100000    0001110111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07645 - 07649

  --0001110111100010    0001110111100011    0001110111100100    0001110111100101    0001110111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07650 - 07654

  --0001110111100111    0001110111101000    0001110111101001    0001110111101010    0001110111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07655 - 07659

  --0001110111101100    0001110111101101    0001110111101110    0001110111101111    0001110111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07660 - 07664

  --0001110111110001    0001110111110010    0001110111110011    0001110111110100    0001110111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07665 - 07669

  --0001110111110110    0001110111110111    0001110111111000    0001110111111001    0001110111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07670 - 07674

  --0001110111111011    0001110111111100    0001110111111101    0001110111111110    0001110111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07675 - 07679

  --0001111000000000    0001111000000001    0001111000000010    0001111000000011    0001111000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07680 - 07684

  --0001111000000101    0001111000000110    0001111000000111    0001111000001000    0001111000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07685 - 07689

  --0001111000001010    0001111000001011    0001111000001100    0001111000001101    0001111000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07690 - 07694

  --0001111000001111    0001111000010000    0001111000010001    0001111000010010    0001111000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07695 - 07699

  --0001111000010100    0001111000010101    0001111000010110    0001111000010111    0001111000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07700 - 07704

  --0001111000011001    0001111000011010    0001111000011011    0001111000011100    0001111000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07705 - 07709

  --0001111000011110    0001111000011111    0001111000100000    0001111000100001    0001111000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07710 - 07714

  --0001111000100011    0001111000100100    0001111000100101    0001111000100110    0001111000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07715 - 07719

  --0001111000101000    0001111000101001    0001111000101010    0001111000101011    0001111000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07720 - 07724

  --0001111000101101    0001111000101110    0001111000101111    0001111000110000    0001111000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07725 - 07729

  --0001111000110010    0001111000110011    0001111000110100    0001111000110101    0001111000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07730 - 07734

  --0001111000110111    0001111000111000    0001111000111001    0001111000111010    0001111000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07735 - 07739

  --0001111000111100    0001111000111101    0001111000111110    0001111000111111    0001111001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07740 - 07744

  --0001111001000001    0001111001000010    0001111001000011    0001111001000100    0001111001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07745 - 07749

  --0001111001000110    0001111001000111    0001111001001000    0001111001001001    0001111001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07750 - 07754

  --0001111001001011    0001111001001100    0001111001001101    0001111001001110    0001111001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07755 - 07759

  --0001111001010000    0001111001010001    0001111001010010    0001111001010011    0001111001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07760 - 07764

  --0001111001010101    0001111001010110    0001111001010111    0001111001011000    0001111001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07765 - 07769

  --0001111001011010    0001111001011011    0001111001011100    0001111001011101    0001111001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07770 - 07774

  --0001111001011111    0001111001100000    0001111001100001    0001111001100010    0001111001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07775 - 07779

  --0001111001100100    0001111001100101    0001111001100110    0001111001100111    0001111001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07780 - 07784

  --0001111001101001    0001111001101010    0001111001101011    0001111001101100    0001111001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07785 - 07789

  --0001111001101110    0001111001101111    0001111001110000    0001111001110001    0001111001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07790 - 07794

  --0001111001110011    0001111001110100    0001111001110101    0001111001110110    0001111001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07795 - 07799

  --0001111001111000    0001111001111001    0001111001111010    0001111001111011    0001111001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07800 - 07804

  --0001111001111101    0001111001111110    0001111001111111    0001111010000000    0001111010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07805 - 07809

  --0001111010000010    0001111010000011    0001111010000100    0001111010000101    0001111010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07810 - 07814

  --0001111010000111    0001111010001000    0001111010001001    0001111010001010    0001111010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07815 - 07819

  --0001111010001100    0001111010001101    0001111010001110    0001111010001111    0001111010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07820 - 07824

  --0001111010010001    0001111010010010    0001111010010011    0001111010010100    0001111010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07825 - 07829

  --0001111010010110    0001111010010111    0001111010011000    0001111010011001    0001111010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07830 - 07834

  --0001111010011011    0001111010011100    0001111010011101    0001111010011110    0001111010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07835 - 07839

  --0001111010100000    0001111010100001    0001111010100010    0001111010100011    0001111010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07840 - 07844

  --0001111010100101    0001111010100110    0001111010100111    0001111010101000    0001111010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07845 - 07849

  --0001111010101010    0001111010101011    0001111010101100    0001111010101101    0001111010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07850 - 07854

  --0001111010101111    0001111010110000    0001111010110001    0001111010110010    0001111010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07855 - 07859

  --0001111010110100    0001111010110101    0001111010110110    0001111010110111    0001111010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07860 - 07864

  --0001111010111001    0001111010111010    0001111010111011    0001111010111100    0001111010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07865 - 07869

  --0001111010111110    0001111010111111    0001111011000000    0001111011000001    0001111011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07870 - 07874

  --0001111011000011    0001111011000100    0001111011000101    0001111011000110    0001111011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07875 - 07879

  --0001111011001000    0001111011001001    0001111011001010    0001111011001011    0001111011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07880 - 07884

  --0001111011001101    0001111011001110    0001111011001111    0001111011010000    0001111011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07885 - 07889

  --0001111011010010    0001111011010011    0001111011010100    0001111011010101    0001111011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07890 - 07894

  --0001111011010111    0001111011011000    0001111011011001    0001111011011010    0001111011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07895 - 07899

  --0001111011011100    0001111011011101    0001111011011110    0001111011011111    0001111011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07900 - 07904

  --0001111011100001    0001111011100010    0001111011100011    0001111011100100    0001111011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07905 - 07909

  --0001111011100110    0001111011100111    0001111011101000    0001111011101001    0001111011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07910 - 07914

  --0001111011101011    0001111011101100    0001111011101101    0001111011101110    0001111011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07915 - 07919

  --0001111011110000    0001111011110001    0001111011110010    0001111011110011    0001111011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07920 - 07924

  --0001111011110101    0001111011110110    0001111011110111    0001111011111000    0001111011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07925 - 07929

  --0001111011111010    0001111011111011    0001111011111100    0001111011111101    0001111011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07930 - 07934

  --0001111011111111    0001111100000000    0001111100000001    0001111100000010    0001111100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07935 - 07939

  --0001111100000100    0001111100000101    0001111100000110    0001111100000111    0001111100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07940 - 07944

  --0001111100001001    0001111100001010    0001111100001011    0001111100001100    0001111100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07945 - 07949

  --0001111100001110    0001111100001111    0001111100010000    0001111100010001    0001111100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07950 - 07954

  --0001111100010011    0001111100010100    0001111100010101    0001111100010110    0001111100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07955 - 07959

  --0001111100011000    0001111100011001    0001111100011010    0001111100011011    0001111100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07960 - 07964

  --0001111100011101    0001111100011110    0001111100011111    0001111100100000    0001111100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07965 - 07969

  --0001111100100010    0001111100100011    0001111100100100    0001111100100101    0001111100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07970 - 07974

  --0001111100100111    0001111100101000    0001111100101001    0001111100101010    0001111100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07975 - 07979

  --0001111100101100    0001111100101101    0001111100101110    0001111100101111    0001111100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07980 - 07984

  --0001111100110001    0001111100110010    0001111100110011    0001111100110100    0001111100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07985 - 07989

  --0001111100110110    0001111100110111    0001111100111000    0001111100111001    0001111100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07990 - 07994

  --0001111100111011    0001111100111100    0001111100111101    0001111100111110    0001111100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 07995 - 07999

  --0001111101000000    0001111101000001    0001111101000010    0001111101000011    0001111101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08000 - 08004

  --0001111101000101    0001111101000110    0001111101000111    0001111101001000    0001111101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08005 - 08009

  --0001111101001010    0001111101001011    0001111101001100    0001111101001101    0001111101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08010 - 08014

  --0001111101001111    0001111101010000    0001111101010001    0001111101010010    0001111101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08015 - 08019

  --0001111101010100    0001111101010101    0001111101010110    0001111101010111    0001111101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08020 - 08024

  --0001111101011001    0001111101011010    0001111101011011    0001111101011100    0001111101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08025 - 08029

  --0001111101011110    0001111101011111    0001111101100000    0001111101100001    0001111101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08030 - 08034

  --0001111101100011    0001111101100100    0001111101100101    0001111101100110    0001111101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08035 - 08039

  --0001111101101000    0001111101101001    0001111101101010    0001111101101011    0001111101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08040 - 08044

  --0001111101101101    0001111101101110    0001111101101111    0001111101110000    0001111101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08045 - 08049

  --0001111101110010    0001111101110011    0001111101110100    0001111101110101    0001111101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08050 - 08054

  --0001111101110111    0001111101111000    0001111101111001    0001111101111010    0001111101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08055 - 08059

  --0001111101111100    0001111101111101    0001111101111110    0001111101111111    0001111110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08060 - 08064

  --0001111110000001    0001111110000010    0001111110000011    0001111110000100    0001111110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08065 - 08069

  --0001111110000110    0001111110000111    0001111110001000    0001111110001001    0001111110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08070 - 08074

  --0001111110001011    0001111110001100    0001111110001101    0001111110001110    0001111110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08075 - 08079

  --0001111110010000    0001111110010001    0001111110010010    0001111110010011    0001111110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08080 - 08084

  --0001111110010101    0001111110010110    0001111110010111    0001111110011000    0001111110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08085 - 08089

  --0001111110011010    0001111110011011    0001111110011100    0001111110011101    0001111110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08090 - 08094

  --0001111110011111    0001111110100000    0001111110100001    0001111110100010    0001111110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08095 - 08099

  --0001111110100100    0001111110100101    0001111110100110    0001111110100111    0001111110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08100 - 08104

  --0001111110101001    0001111110101010    0001111110101011    0001111110101100    0001111110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08105 - 08109

  --0001111110101110    0001111110101111    0001111110110000    0001111110110001    0001111110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08110 - 08114

  --0001111110110011    0001111110110100    0001111110110101    0001111110110110    0001111110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08115 - 08119

  --0001111110111000    0001111110111001    0001111110111010    0001111110111011    0001111110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08120 - 08124

  --0001111110111101    0001111110111110    0001111110111111    0001111111000000    0001111111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08125 - 08129

  --0001111111000010    0001111111000011    0001111111000100    0001111111000101    0001111111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08130 - 08134

  --0001111111000111    0001111111001000    0001111111001001    0001111111001010    0001111111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08135 - 08139

  --0001111111001100    0001111111001101    0001111111001110    0001111111001111    0001111111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08140 - 08144

  --0001111111010001    0001111111010010    0001111111010011    0001111111010100    0001111111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08145 - 08149

  --0001111111010110    0001111111010111    0001111111011000    0001111111011001    0001111111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08150 - 08154

  --0001111111011011    0001111111011100    0001111111011101    0001111111011110    0001111111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08155 - 08159

  --0001111111100000    0001111111100001    0001111111100010    0001111111100011    0001111111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08160 - 08164

  --0001111111100101    0001111111100110    0001111111100111    0001111111101000    0001111111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08165 - 08169

  --0001111111101010    0001111111101011    0001111111101100    0001111111101101    0001111111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08170 - 08174

  --0001111111101111    0001111111110000    0001111111110001    0001111111110010    0001111111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08175 - 08179

  --0001111111110100    0001111111110101    0001111111110110    0001111111110111    0001111111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08180 - 08184

  --0001111111111001    0001111111111010    0001111111111011    0001111111111100    0001111111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08185 - 08189

  --0001111111111110    0001111111111111    0010000000000000    0010000000000001    0010000000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08190 - 08194

  --0010000000000011    0010000000000100    0010000000000101    0010000000000110    0010000000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08195 - 08199

  --0010000000001000    0010000000001001    0010000000001010    0010000000001011    0010000000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08200 - 08204

  --0010000000001101    0010000000001110    0010000000001111    0010000000010000    0010000000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08205 - 08209

  --0010000000010010    0010000000010011    0010000000010100    0010000000010101    0010000000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08210 - 08214

  --0010000000010111    0010000000011000    0010000000011001    0010000000011010    0010000000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08215 - 08219

  --0010000000011100    0010000000011101    0010000000011110    0010000000011111    0010000000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08220 - 08224

  --0010000000100001    0010000000100010    0010000000100011    0010000000100100    0010000000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08225 - 08229

  --0010000000100110    0010000000100111    0010000000101000    0010000000101001    0010000000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08230 - 08234

  --0010000000101011    0010000000101100    0010000000101101    0010000000101110    0010000000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08235 - 08239

  --0010000000110000    0010000000110001    0010000000110010    0010000000110011    0010000000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08240 - 08244

  --0010000000110101    0010000000110110    0010000000110111    0010000000111000    0010000000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08245 - 08249

  --0010000000111010    0010000000111011    0010000000111100    0010000000111101    0010000000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08250 - 08254

  --0010000000111111    0010000001000000    0010000001000001    0010000001000010    0010000001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08255 - 08259

  --0010000001000100    0010000001000101    0010000001000110    0010000001000111    0010000001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08260 - 08264

  --0010000001001001    0010000001001010    0010000001001011    0010000001001100    0010000001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08265 - 08269

  --0010000001001110    0010000001001111    0010000001010000    0010000001010001    0010000001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08270 - 08274

  --0010000001010011    0010000001010100    0010000001010101    0010000001010110    0010000001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08275 - 08279

  --0010000001011000    0010000001011001    0010000001011010    0010000001011011    0010000001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08280 - 08284

  --0010000001011101    0010000001011110    0010000001011111    0010000001100000    0010000001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08285 - 08289

  --0010000001100010    0010000001100011    0010000001100100    0010000001100101    0010000001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08290 - 08294

  --0010000001100111    0010000001101000    0010000001101001    0010000001101010    0010000001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08295 - 08299

  --0010000001101100    0010000001101101    0010000001101110    0010000001101111    0010000001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08300 - 08304

  --0010000001110001    0010000001110010    0010000001110011    0010000001110100    0010000001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08305 - 08309

  --0010000001110110    0010000001110111    0010000001111000    0010000001111001    0010000001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08310 - 08314

  --0010000001111011    0010000001111100    0010000001111101    0010000001111110    0010000001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08315 - 08319

  --0010000010000000    0010000010000001    0010000010000010    0010000010000011    0010000010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08320 - 08324

  --0010000010000101    0010000010000110    0010000010000111    0010000010001000    0010000010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08325 - 08329

  --0010000010001010    0010000010001011    0010000010001100    0010000010001101    0010000010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08330 - 08334

  --0010000010001111    0010000010010000    0010000010010001    0010000010010010    0010000010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08335 - 08339

  --0010000010010100    0010000010010101    0010000010010110    0010000010010111    0010000010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08340 - 08344

  --0010000010011001    0010000010011010    0010000010011011    0010000010011100    0010000010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08345 - 08349

  --0010000010011110    0010000010011111    0010000010100000    0010000010100001    0010000010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08350 - 08354

  --0010000010100011    0010000010100100    0010000010100101    0010000010100110    0010000010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08355 - 08359

  --0010000010101000    0010000010101001    0010000010101010    0010000010101011    0010000010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08360 - 08364

  --0010000010101101    0010000010101110    0010000010101111    0010000010110000    0010000010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08365 - 08369

  --0010000010110010    0010000010110011    0010000010110100    0010000010110101    0010000010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08370 - 08374

  --0010000010110111    0010000010111000    0010000010111001    0010000010111010    0010000010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08375 - 08379

  --0010000010111100    0010000010111101    0010000010111110    0010000010111111    0010000011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08380 - 08384

  --0010000011000001    0010000011000010    0010000011000011    0010000011000100    0010000011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08385 - 08389

  --0010000011000110    0010000011000111    0010000011001000    0010000011001001    0010000011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08390 - 08394

  --0010000011001011    0010000011001100    0010000011001101    0010000011001110    0010000011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08395 - 08399

  --0010000011010000    0010000011010001    0010000011010010    0010000011010011    0010000011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08400 - 08404

  --0010000011010101    0010000011010110    0010000011010111    0010000011011000    0010000011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08405 - 08409

  --0010000011011010    0010000011011011    0010000011011100    0010000011011101    0010000011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08410 - 08414

  --0010000011011111    0010000011100000    0010000011100001    0010000011100010    0010000011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08415 - 08419

  --0010000011100100    0010000011100101    0010000011100110    0010000011100111    0010000011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08420 - 08424

  --0010000011101001    0010000011101010    0010000011101011    0010000011101100    0010000011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08425 - 08429

  --0010000011101110    0010000011101111    0010000011110000    0010000011110001    0010000011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08430 - 08434

  --0010000011110011    0010000011110100    0010000011110101    0010000011110110    0010000011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08435 - 08439

  --0010000011111000    0010000011111001    0010000011111010    0010000011111011    0010000011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08440 - 08444

  --0010000011111101    0010000011111110    0010000011111111    0010000100000000    0010000100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08445 - 08449

  --0010000100000010    0010000100000011    0010000100000100    0010000100000101    0010000100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08450 - 08454

  --0010000100000111    0010000100001000    0010000100001001    0010000100001010    0010000100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08455 - 08459

  --0010000100001100    0010000100001101    0010000100001110    0010000100001111    0010000100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08460 - 08464

  --0010000100010001    0010000100010010    0010000100010011    0010000100010100    0010000100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08465 - 08469

  --0010000100010110    0010000100010111    0010000100011000    0010000100011001    0010000100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08470 - 08474

  --0010000100011011    0010000100011100    0010000100011101    0010000100011110    0010000100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08475 - 08479

  --0010000100100000    0010000100100001    0010000100100010    0010000100100011    0010000100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08480 - 08484

  --0010000100100101    0010000100100110    0010000100100111    0010000100101000    0010000100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08485 - 08489

  --0010000100101010    0010000100101011    0010000100101100    0010000100101101    0010000100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08490 - 08494

  --0010000100101111    0010000100110000    0010000100110001    0010000100110010    0010000100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08495 - 08499

  --0010000100110100    0010000100110101    0010000100110110    0010000100110111    0010000100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08500 - 08504

  --0010000100111001    0010000100111010    0010000100111011    0010000100111100    0010000100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08505 - 08509

  --0010000100111110    0010000100111111    0010000101000000    0010000101000001    0010000101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08510 - 08514

  --0010000101000011    0010000101000100    0010000101000101    0010000101000110    0010000101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08515 - 08519

  --0010000101001000    0010000101001001    0010000101001010    0010000101001011    0010000101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08520 - 08524

  --0010000101001101    0010000101001110    0010000101001111    0010000101010000    0010000101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08525 - 08529

  --0010000101010010    0010000101010011    0010000101010100    0010000101010101    0010000101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08530 - 08534

  --0010000101010111    0010000101011000    0010000101011001    0010000101011010    0010000101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08535 - 08539

  --0010000101011100    0010000101011101    0010000101011110    0010000101011111    0010000101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08540 - 08544

  --0010000101100001    0010000101100010    0010000101100011    0010000101100100    0010000101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08545 - 08549

  --0010000101100110    0010000101100111    0010000101101000    0010000101101001    0010000101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08550 - 08554

  --0010000101101011    0010000101101100    0010000101101101    0010000101101110    0010000101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08555 - 08559

  --0010000101110000    0010000101110001    0010000101110010    0010000101110011    0010000101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08560 - 08564

  --0010000101110101    0010000101110110    0010000101110111    0010000101111000    0010000101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08565 - 08569

  --0010000101111010    0010000101111011    0010000101111100    0010000101111101    0010000101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08570 - 08574

  --0010000101111111    0010000110000000    0010000110000001    0010000110000010    0010000110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08575 - 08579

  --0010000110000100    0010000110000101    0010000110000110    0010000110000111    0010000110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08580 - 08584

  --0010000110001001    0010000110001010    0010000110001011    0010000110001100    0010000110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08585 - 08589

  --0010000110001110    0010000110001111    0010000110010000    0010000110010001    0010000110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08590 - 08594

  --0010000110010011    0010000110010100    0010000110010101    0010000110010110    0010000110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08595 - 08599

  --0010000110011000    0010000110011001    0010000110011010    0010000110011011    0010000110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08600 - 08604

  --0010000110011101    0010000110011110    0010000110011111    0010000110100000    0010000110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08605 - 08609

  --0010000110100010    0010000110100011    0010000110100100    0010000110100101    0010000110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08610 - 08614

  --0010000110100111    0010000110101000    0010000110101001    0010000110101010    0010000110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08615 - 08619

  --0010000110101100    0010000110101101    0010000110101110    0010000110101111    0010000110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08620 - 08624

  --0010000110110001    0010000110110010    0010000110110011    0010000110110100    0010000110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08625 - 08629

  --0010000110110110    0010000110110111    0010000110111000    0010000110111001    0010000110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08630 - 08634

  --0010000110111011    0010000110111100    0010000110111101    0010000110111110    0010000110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08635 - 08639

  --0010000111000000    0010000111000001    0010000111000010    0010000111000011    0010000111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08640 - 08644

  --0010000111000101    0010000111000110    0010000111000111    0010000111001000    0010000111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08645 - 08649

  --0010000111001010    0010000111001011    0010000111001100    0010000111001101    0010000111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08650 - 08654

  --0010000111001111    0010000111010000    0010000111010001    0010000111010010    0010000111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08655 - 08659

  --0010000111010100    0010000111010101    0010000111010110    0010000111010111    0010000111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08660 - 08664

  --0010000111011001    0010000111011010    0010000111011011    0010000111011100    0010000111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08665 - 08669

  --0010000111011110    0010000111011111    0010000111100000    0010000111100001    0010000111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08670 - 08674

  --0010000111100011    0010000111100100    0010000111100101    0010000111100110    0010000111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08675 - 08679

  --0010000111101000    0010000111101001    0010000111101010    0010000111101011    0010000111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08680 - 08684

  --0010000111101101    0010000111101110    0010000111101111    0010000111110000    0010000111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08685 - 08689

  --0010000111110010    0010000111110011    0010000111110100    0010000111110101    0010000111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08690 - 08694

  --0010000111110111    0010000111111000    0010000111111001    0010000111111010    0010000111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08695 - 08699

  --0010000111111100    0010000111111101    0010000111111110    0010000111111111    0010001000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08700 - 08704

  --0010001000000001    0010001000000010    0010001000000011    0010001000000100    0010001000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08705 - 08709

  --0010001000000110    0010001000000111    0010001000001000    0010001000001001    0010001000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08710 - 08714

  --0010001000001011    0010001000001100    0010001000001101    0010001000001110    0010001000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08715 - 08719

  --0010001000010000    0010001000010001    0010001000010010    0010001000010011    0010001000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08720 - 08724

  --0010001000010101    0010001000010110    0010001000010111    0010001000011000    0010001000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08725 - 08729

  --0010001000011010    0010001000011011    0010001000011100    0010001000011101    0010001000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08730 - 08734

  --0010001000011111    0010001000100000    0010001000100001    0010001000100010    0010001000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08735 - 08739

  --0010001000100100    0010001000100101    0010001000100110    0010001000100111    0010001000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08740 - 08744

  --0010001000101001    0010001000101010    0010001000101011    0010001000101100    0010001000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08745 - 08749

  --0010001000101110    0010001000101111    0010001000110000    0010001000110001    0010001000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08750 - 08754

  --0010001000110011    0010001000110100    0010001000110101    0010001000110110    0010001000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08755 - 08759

  --0010001000111000    0010001000111001    0010001000111010    0010001000111011    0010001000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08760 - 08764

  --0010001000111101    0010001000111110    0010001000111111    0010001001000000    0010001001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08765 - 08769

  --0010001001000010    0010001001000011    0010001001000100    0010001001000101    0010001001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08770 - 08774

  --0010001001000111    0010001001001000    0010001001001001    0010001001001010    0010001001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08775 - 08779

  --0010001001001100    0010001001001101    0010001001001110    0010001001001111    0010001001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08780 - 08784

  --0010001001010001    0010001001010010    0010001001010011    0010001001010100    0010001001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08785 - 08789

  --0010001001010110    0010001001010111    0010001001011000    0010001001011001    0010001001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08790 - 08794

  --0010001001011011    0010001001011100    0010001001011101    0010001001011110    0010001001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08795 - 08799

  --0010001001100000    0010001001100001    0010001001100010    0010001001100011    0010001001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08800 - 08804

  --0010001001100101    0010001001100110    0010001001100111    0010001001101000    0010001001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08805 - 08809

  --0010001001101010    0010001001101011    0010001001101100    0010001001101101    0010001001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08810 - 08814

  --0010001001101111    0010001001110000    0010001001110001    0010001001110010    0010001001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08815 - 08819

  --0010001001110100    0010001001110101    0010001001110110    0010001001110111    0010001001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08820 - 08824

  --0010001001111001    0010001001111010    0010001001111011    0010001001111100    0010001001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08825 - 08829

  --0010001001111110    0010001001111111    0010001010000000    0010001010000001    0010001010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08830 - 08834

  --0010001010000011    0010001010000100    0010001010000101    0010001010000110    0010001010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08835 - 08839

  --0010001010001000    0010001010001001    0010001010001010    0010001010001011    0010001010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08840 - 08844

  --0010001010001101    0010001010001110    0010001010001111    0010001010010000    0010001010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08845 - 08849

  --0010001010010010    0010001010010011    0010001010010100    0010001010010101    0010001010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08850 - 08854

  --0010001010010111    0010001010011000    0010001010011001    0010001010011010    0010001010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08855 - 08859

  --0010001010011100    0010001010011101    0010001010011110    0010001010011111    0010001010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08860 - 08864

  --0010001010100001    0010001010100010    0010001010100011    0010001010100100    0010001010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08865 - 08869

  --0010001010100110    0010001010100111    0010001010101000    0010001010101001    0010001010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08870 - 08874

  --0010001010101011    0010001010101100    0010001010101101    0010001010101110    0010001010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08875 - 08879

  --0010001010110000    0010001010110001    0010001010110010    0010001010110011    0010001010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08880 - 08884

  --0010001010110101    0010001010110110    0010001010110111    0010001010111000    0010001010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08885 - 08889

  --0010001010111010    0010001010111011    0010001010111100    0010001010111101    0010001010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08890 - 08894

  --0010001010111111    0010001011000000    0010001011000001    0010001011000010    0010001011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08895 - 08899

  --0010001011000100    0010001011000101    0010001011000110    0010001011000111    0010001011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08900 - 08904

  --0010001011001001    0010001011001010    0010001011001011    0010001011001100    0010001011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08905 - 08909

  --0010001011001110    0010001011001111    0010001011010000    0010001011010001    0010001011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08910 - 08914

  --0010001011010011    0010001011010100    0010001011010101    0010001011010110    0010001011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08915 - 08919

  --0010001011011000    0010001011011001    0010001011011010    0010001011011011    0010001011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08920 - 08924

  --0010001011011101    0010001011011110    0010001011011111    0010001011100000    0010001011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08925 - 08929

  --0010001011100010    0010001011100011    0010001011100100    0010001011100101    0010001011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08930 - 08934

  --0010001011100111    0010001011101000    0010001011101001    0010001011101010    0010001011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08935 - 08939

  --0010001011101100    0010001011101101    0010001011101110    0010001011101111    0010001011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08940 - 08944

  --0010001011110001    0010001011110010    0010001011110011    0010001011110100    0010001011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08945 - 08949

  --0010001011110110    0010001011110111    0010001011111000    0010001011111001    0010001011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08950 - 08954

  --0010001011111011    0010001011111100    0010001011111101    0010001011111110    0010001011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08955 - 08959

  --0010001100000000    0010001100000001    0010001100000010    0010001100000011    0010001100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08960 - 08964

  --0010001100000101    0010001100000110    0010001100000111    0010001100001000    0010001100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08965 - 08969

  --0010001100001010    0010001100001011    0010001100001100    0010001100001101    0010001100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08970 - 08974

  --0010001100001111    0010001100010000    0010001100010001    0010001100010010    0010001100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08975 - 08979

  --0010001100010100    0010001100010101    0010001100010110    0010001100010111    0010001100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08980 - 08984

  --0010001100011001    0010001100011010    0010001100011011    0010001100011100    0010001100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08985 - 08989

  --0010001100011110    0010001100011111    0010001100100000    0010001100100001    0010001100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08990 - 08994

  --0010001100100011    0010001100100100    0010001100100101    0010001100100110    0010001100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 08995 - 08999

  --0010001100101000    0010001100101001    0010001100101010    0010001100101011    0010001100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09000 - 09004

  --0010001100101101    0010001100101110    0010001100101111    0010001100110000    0010001100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09005 - 09009

  --0010001100110010    0010001100110011    0010001100110100    0010001100110101    0010001100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09010 - 09014

  --0010001100110111    0010001100111000    0010001100111001    0010001100111010    0010001100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09015 - 09019

  --0010001100111100    0010001100111101    0010001100111110    0010001100111111    0010001101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09020 - 09024

  --0010001101000001    0010001101000010    0010001101000011    0010001101000100    0010001101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09025 - 09029

  --0010001101000110    0010001101000111    0010001101001000    0010001101001001    0010001101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09030 - 09034

  --0010001101001011    0010001101001100    0010001101001101    0010001101001110    0010001101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09035 - 09039

  --0010001101010000    0010001101010001    0010001101010010    0010001101010011    0010001101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09040 - 09044

  --0010001101010101    0010001101010110    0010001101010111    0010001101011000    0010001101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09045 - 09049

  --0010001101011010    0010001101011011    0010001101011100    0010001101011101    0010001101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09050 - 09054

  --0010001101011111    0010001101100000    0010001101100001    0010001101100010    0010001101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09055 - 09059

  --0010001101100100    0010001101100101    0010001101100110    0010001101100111    0010001101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09060 - 09064

  --0010001101101001    0010001101101010    0010001101101011    0010001101101100    0010001101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09065 - 09069

  --0010001101101110    0010001101101111    0010001101110000    0010001101110001    0010001101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09070 - 09074

  --0010001101110011    0010001101110100    0010001101110101    0010001101110110    0010001101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09075 - 09079

  --0010001101111000    0010001101111001    0010001101111010    0010001101111011    0010001101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09080 - 09084

  --0010001101111101    0010001101111110    0010001101111111    0010001110000000    0010001110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09085 - 09089

  --0010001110000010    0010001110000011    0010001110000100    0010001110000101    0010001110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09090 - 09094

  --0010001110000111    0010001110001000    0010001110001001    0010001110001010    0010001110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09095 - 09099

  --0010001110001100    0010001110001101    0010001110001110    0010001110001111    0010001110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09100 - 09104

  --0010001110010001    0010001110010010    0010001110010011    0010001110010100    0010001110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09105 - 09109

  --0010001110010110    0010001110010111    0010001110011000    0010001110011001    0010001110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09110 - 09114

  --0010001110011011    0010001110011100    0010001110011101    0010001110011110    0010001110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09115 - 09119

  --0010001110100000    0010001110100001    0010001110100010    0010001110100011    0010001110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09120 - 09124

  --0010001110100101    0010001110100110    0010001110100111    0010001110101000    0010001110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09125 - 09129

  --0010001110101010    0010001110101011    0010001110101100    0010001110101101    0010001110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09130 - 09134

  --0010001110101111    0010001110110000    0010001110110001    0010001110110010    0010001110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09135 - 09139

  --0010001110110100    0010001110110101    0010001110110110    0010001110110111    0010001110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09140 - 09144

  --0010001110111001    0010001110111010    0010001110111011    0010001110111100    0010001110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09145 - 09149

  --0010001110111110    0010001110111111    0010001111000000    0010001111000001    0010001111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09150 - 09154

  --0010001111000011    0010001111000100    0010001111000101    0010001111000110    0010001111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09155 - 09159

  --0010001111001000    0010001111001001    0010001111001010    0010001111001011    0010001111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09160 - 09164

  --0010001111001101    0010001111001110    0010001111001111    0010001111010000    0010001111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09165 - 09169

  --0010001111010010    0010001111010011    0010001111010100    0010001111010101    0010001111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09170 - 09174

  --0010001111010111    0010001111011000    0010001111011001    0010001111011010    0010001111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09175 - 09179

  --0010001111011100    0010001111011101    0010001111011110    0010001111011111    0010001111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09180 - 09184

  --0010001111100001    0010001111100010    0010001111100011    0010001111100100    0010001111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09185 - 09189

  --0010001111100110    0010001111100111    0010001111101000    0010001111101001    0010001111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09190 - 09194

  --0010001111101011    0010001111101100    0010001111101101    0010001111101110    0010001111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09195 - 09199

  --0010001111110000    0010001111110001    0010001111110010    0010001111110011    0010001111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09200 - 09204

  --0010001111110101    0010001111110110    0010001111110111    0010001111111000    0010001111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09205 - 09209

  --0010001111111010    0010001111111011    0010001111111100    0010001111111101    0010001111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09210 - 09214

  --0010001111111111    0010010000000000    0010010000000001    0010010000000010    0010010000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09215 - 09219

  --0010010000000100    0010010000000101    0010010000000110    0010010000000111    0010010000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09220 - 09224

  --0010010000001001    0010010000001010    0010010000001011    0010010000001100    0010010000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09225 - 09229

  --0010010000001110    0010010000001111    0010010000010000    0010010000010001    0010010000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09230 - 09234

  --0010010000010011    0010010000010100    0010010000010101    0010010000010110    0010010000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09235 - 09239

  --0010010000011000    0010010000011001    0010010000011010    0010010000011011    0010010000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09240 - 09244

  --0010010000011101    0010010000011110    0010010000011111    0010010000100000    0010010000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09245 - 09249

  --0010010000100010    0010010000100011    0010010000100100    0010010000100101    0010010000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09250 - 09254

  --0010010000100111    0010010000101000    0010010000101001    0010010000101010    0010010000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09255 - 09259

  --0010010000101100    0010010000101101    0010010000101110    0010010000101111    0010010000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09260 - 09264

  --0010010000110001    0010010000110010    0010010000110011    0010010000110100    0010010000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09265 - 09269

  --0010010000110110    0010010000110111    0010010000111000    0010010000111001    0010010000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09270 - 09274

  --0010010000111011    0010010000111100    0010010000111101    0010010000111110    0010010000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09275 - 09279

  --0010010001000000    0010010001000001    0010010001000010    0010010001000011    0010010001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09280 - 09284

  --0010010001000101    0010010001000110    0010010001000111    0010010001001000    0010010001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09285 - 09289

  --0010010001001010    0010010001001011    0010010001001100    0010010001001101    0010010001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09290 - 09294

  --0010010001001111    0010010001010000    0010010001010001    0010010001010010    0010010001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09295 - 09299

  --0010010001010100    0010010001010101    0010010001010110    0010010001010111    0010010001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09300 - 09304

  --0010010001011001    0010010001011010    0010010001011011    0010010001011100    0010010001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09305 - 09309

  --0010010001011110    0010010001011111    0010010001100000    0010010001100001    0010010001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09310 - 09314

  --0010010001100011    0010010001100100    0010010001100101    0010010001100110    0010010001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09315 - 09319

  --0010010001101000    0010010001101001    0010010001101010    0010010001101011    0010010001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09320 - 09324

  --0010010001101101    0010010001101110    0010010001101111    0010010001110000    0010010001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09325 - 09329

  --0010010001110010    0010010001110011    0010010001110100    0010010001110101    0010010001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09330 - 09334

  --0010010001110111    0010010001111000    0010010001111001    0010010001111010    0010010001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09335 - 09339

  --0010010001111100    0010010001111101    0010010001111110    0010010001111111    0010010010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09340 - 09344

  --0010010010000001    0010010010000010    0010010010000011    0010010010000100    0010010010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09345 - 09349

  --0010010010000110    0010010010000111    0010010010001000    0010010010001001    0010010010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09350 - 09354

  --0010010010001011    0010010010001100    0010010010001101    0010010010001110    0010010010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09355 - 09359

  --0010010010010000    0010010010010001    0010010010010010    0010010010010011    0010010010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09360 - 09364

  --0010010010010101    0010010010010110    0010010010010111    0010010010011000    0010010010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09365 - 09369

  --0010010010011010    0010010010011011    0010010010011100    0010010010011101    0010010010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09370 - 09374

  --0010010010011111    0010010010100000    0010010010100001    0010010010100010    0010010010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09375 - 09379

  --0010010010100100    0010010010100101    0010010010100110    0010010010100111    0010010010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09380 - 09384

  --0010010010101001    0010010010101010    0010010010101011    0010010010101100    0010010010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09385 - 09389

  --0010010010101110    0010010010101111    0010010010110000    0010010010110001    0010010010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09390 - 09394

  --0010010010110011    0010010010110100    0010010010110101    0010010010110110    0010010010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09395 - 09399

  --0010010010111000    0010010010111001    0010010010111010    0010010010111011    0010010010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09400 - 09404

  --0010010010111101    0010010010111110    0010010010111111    0010010011000000    0010010011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09405 - 09409

  --0010010011000010    0010010011000011    0010010011000100    0010010011000101    0010010011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09410 - 09414

  --0010010011000111    0010010011001000    0010010011001001    0010010011001010    0010010011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09415 - 09419

  --0010010011001100    0010010011001101    0010010011001110    0010010011001111    0010010011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09420 - 09424

  --0010010011010001    0010010011010010    0010010011010011    0010010011010100    0010010011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09425 - 09429

  --0010010011010110    0010010011010111    0010010011011000    0010010011011001    0010010011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09430 - 09434

  --0010010011011011    0010010011011100    0010010011011101    0010010011011110    0010010011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09435 - 09439

  --0010010011100000    0010010011100001    0010010011100010    0010010011100011    0010010011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09440 - 09444

  --0010010011100101    0010010011100110    0010010011100111    0010010011101000    0010010011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09445 - 09449

  --0010010011101010    0010010011101011    0010010011101100    0010010011101101    0010010011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09450 - 09454

  --0010010011101111    0010010011110000    0010010011110001    0010010011110010    0010010011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09455 - 09459

  --0010010011110100    0010010011110101    0010010011110110    0010010011110111    0010010011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09460 - 09464

  --0010010011111001    0010010011111010    0010010011111011    0010010011111100    0010010011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09465 - 09469

  --0010010011111110    0010010011111111    0010010100000000    0010010100000001    0010010100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09470 - 09474

  --0010010100000011    0010010100000100    0010010100000101    0010010100000110    0010010100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09475 - 09479

  --0010010100001000    0010010100001001    0010010100001010    0010010100001011    0010010100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09480 - 09484

  --0010010100001101    0010010100001110    0010010100001111    0010010100010000    0010010100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09485 - 09489

  --0010010100010010    0010010100010011    0010010100010100    0010010100010101    0010010100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09490 - 09494

  --0010010100010111    0010010100011000    0010010100011001    0010010100011010    0010010100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09495 - 09499

  --0010010100011100    0010010100011101    0010010100011110    0010010100011111    0010010100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09500 - 09504

  --0010010100100001    0010010100100010    0010010100100011    0010010100100100    0010010100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09505 - 09509

  --0010010100100110    0010010100100111    0010010100101000    0010010100101001    0010010100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09510 - 09514

  --0010010100101011    0010010100101100    0010010100101101    0010010100101110    0010010100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09515 - 09519

  --0010010100110000    0010010100110001    0010010100110010    0010010100110011    0010010100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09520 - 09524

  --0010010100110101    0010010100110110    0010010100110111    0010010100111000    0010010100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09525 - 09529

  --0010010100111010    0010010100111011    0010010100111100    0010010100111101    0010010100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09530 - 09534

  --0010010100111111    0010010101000000    0010010101000001    0010010101000010    0010010101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09535 - 09539

  --0010010101000100    0010010101000101    0010010101000110    0010010101000111    0010010101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09540 - 09544

  --0010010101001001    0010010101001010    0010010101001011    0010010101001100    0010010101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09545 - 09549

  --0010010101001110    0010010101001111    0010010101010000    0010010101010001    0010010101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09550 - 09554

  --0010010101010011    0010010101010100    0010010101010101    0010010101010110    0010010101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09555 - 09559

  --0010010101011000    0010010101011001    0010010101011010    0010010101011011    0010010101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09560 - 09564

  --0010010101011101    0010010101011110    0010010101011111    0010010101100000    0010010101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09565 - 09569

  --0010010101100010    0010010101100011    0010010101100100    0010010101100101    0010010101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09570 - 09574

  --0010010101100111    0010010101101000    0010010101101001    0010010101101010    0010010101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09575 - 09579

  --0010010101101100    0010010101101101    0010010101101110    0010010101101111    0010010101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09580 - 09584

  --0010010101110001    0010010101110010    0010010101110011    0010010101110100    0010010101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09585 - 09589

  --0010010101110110    0010010101110111    0010010101111000    0010010101111001    0010010101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09590 - 09594

  --0010010101111011    0010010101111100    0010010101111101    0010010101111110    0010010101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09595 - 09599

  --0010010110000000    0010010110000001    0010010110000010    0010010110000011    0010010110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09600 - 09604

  --0010010110000101    0010010110000110    0010010110000111    0010010110001000    0010010110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09605 - 09609

  --0010010110001010    0010010110001011    0010010110001100    0010010110001101    0010010110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09610 - 09614

  --0010010110001111    0010010110010000    0010010110010001    0010010110010010    0010010110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09615 - 09619

  --0010010110010100    0010010110010101    0010010110010110    0010010110010111    0010010110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09620 - 09624

  --0010010110011001    0010010110011010    0010010110011011    0010010110011100    0010010110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09625 - 09629

  --0010010110011110    0010010110011111    0010010110100000    0010010110100001    0010010110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09630 - 09634

  --0010010110100011    0010010110100100    0010010110100101    0010010110100110    0010010110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09635 - 09639

  --0010010110101000    0010010110101001    0010010110101010    0010010110101011    0010010110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09640 - 09644

  --0010010110101101    0010010110101110    0010010110101111    0010010110110000    0010010110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09645 - 09649

  --0010010110110010    0010010110110011    0010010110110100    0010010110110101    0010010110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09650 - 09654

  --0010010110110111    0010010110111000    0010010110111001    0010010110111010    0010010110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09655 - 09659

  --0010010110111100    0010010110111101    0010010110111110    0010010110111111    0010010111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09660 - 09664

  --0010010111000001    0010010111000010    0010010111000011    0010010111000100    0010010111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09665 - 09669

  --0010010111000110    0010010111000111    0010010111001000    0010010111001001    0010010111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09670 - 09674

  --0010010111001011    0010010111001100    0010010111001101    0010010111001110    0010010111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09675 - 09679

  --0010010111010000    0010010111010001    0010010111010010    0010010111010011    0010010111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09680 - 09684

  --0010010111010101    0010010111010110    0010010111010111    0010010111011000    0010010111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09685 - 09689

  --0010010111011010    0010010111011011    0010010111011100    0010010111011101    0010010111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09690 - 09694

  --0010010111011111    0010010111100000    0010010111100001    0010010111100010    0010010111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09695 - 09699

  --0010010111100100    0010010111100101    0010010111100110    0010010111100111    0010010111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09700 - 09704

  --0010010111101001    0010010111101010    0010010111101011    0010010111101100    0010010111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09705 - 09709

  --0010010111101110    0010010111101111    0010010111110000    0010010111110001    0010010111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09710 - 09714

  --0010010111110011    0010010111110100    0010010111110101    0010010111110110    0010010111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09715 - 09719

  --0010010111111000    0010010111111001    0010010111111010    0010010111111011    0010010111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09720 - 09724

  --0010010111111101    0010010111111110    0010010111111111    0010011000000000    0010011000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09725 - 09729

  --0010011000000010    0010011000000011    0010011000000100    0010011000000101    0010011000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09730 - 09734

  --0010011000000111    0010011000001000    0010011000001001    0010011000001010    0010011000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09735 - 09739

  --0010011000001100    0010011000001101    0010011000001110    0010011000001111    0010011000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09740 - 09744

  --0010011000010001    0010011000010010    0010011000010011    0010011000010100    0010011000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09745 - 09749

  --0010011000010110    0010011000010111    0010011000011000    0010011000011001    0010011000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09750 - 09754

  --0010011000011011    0010011000011100    0010011000011101    0010011000011110    0010011000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09755 - 09759

  --0010011000100000    0010011000100001    0010011000100010    0010011000100011    0010011000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09760 - 09764

  --0010011000100101    0010011000100110    0010011000100111    0010011000101000    0010011000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09765 - 09769

  --0010011000101010    0010011000101011    0010011000101100    0010011000101101    0010011000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09770 - 09774

  --0010011000101111    0010011000110000    0010011000110001    0010011000110010    0010011000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09775 - 09779

  --0010011000110100    0010011000110101    0010011000110110    0010011000110111    0010011000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09780 - 09784

  --0010011000111001    0010011000111010    0010011000111011    0010011000111100    0010011000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09785 - 09789

  --0010011000111110    0010011000111111    0010011001000000    0010011001000001    0010011001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09790 - 09794

  --0010011001000011    0010011001000100    0010011001000101    0010011001000110    0010011001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09795 - 09799

  --0010011001001000    0010011001001001    0010011001001010    0010011001001011    0010011001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09800 - 09804

  --0010011001001101    0010011001001110    0010011001001111    0010011001010000    0010011001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09805 - 09809

  --0010011001010010    0010011001010011    0010011001010100    0010011001010101    0010011001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09810 - 09814

  --0010011001010111    0010011001011000    0010011001011001    0010011001011010    0010011001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09815 - 09819

  --0010011001011100    0010011001011101    0010011001011110    0010011001011111    0010011001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09820 - 09824

  --0010011001100001    0010011001100010    0010011001100011    0010011001100100    0010011001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09825 - 09829

  --0010011001100110    0010011001100111    0010011001101000    0010011001101001    0010011001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09830 - 09834

  --0010011001101011    0010011001101100    0010011001101101    0010011001101110    0010011001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09835 - 09839

  --0010011001110000    0010011001110001    0010011001110010    0010011001110011    0010011001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09840 - 09844

  --0010011001110101    0010011001110110    0010011001110111    0010011001111000    0010011001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09845 - 09849

  --0010011001111010    0010011001111011    0010011001111100    0010011001111101    0010011001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09850 - 09854

  --0010011001111111    0010011010000000    0010011010000001    0010011010000010    0010011010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09855 - 09859

  --0010011010000100    0010011010000101    0010011010000110    0010011010000111    0010011010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09860 - 09864

  --0010011010001001    0010011010001010    0010011010001011    0010011010001100    0010011010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09865 - 09869

  --0010011010001110    0010011010001111    0010011010010000    0010011010010001    0010011010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09870 - 09874

  --0010011010010011    0010011010010100    0010011010010101    0010011010010110    0010011010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09875 - 09879

  --0010011010011000    0010011010011001    0010011010011010    0010011010011011    0010011010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09880 - 09884

  --0010011010011101    0010011010011110    0010011010011111    0010011010100000    0010011010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09885 - 09889

  --0010011010100010    0010011010100011    0010011010100100    0010011010100101    0010011010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09890 - 09894

  --0010011010100111    0010011010101000    0010011010101001    0010011010101010    0010011010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09895 - 09899

  --0010011010101100    0010011010101101    0010011010101110    0010011010101111    0010011010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09900 - 09904

  --0010011010110001    0010011010110010    0010011010110011    0010011010110100    0010011010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09905 - 09909

  --0010011010110110    0010011010110111    0010011010111000    0010011010111001    0010011010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09910 - 09914

  --0010011010111011    0010011010111100    0010011010111101    0010011010111110    0010011010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09915 - 09919

  --0010011011000000    0010011011000001    0010011011000010    0010011011000011    0010011011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09920 - 09924

  --0010011011000101    0010011011000110    0010011011000111    0010011011001000    0010011011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09925 - 09929

  --0010011011001010    0010011011001011    0010011011001100    0010011011001101    0010011011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09930 - 09934

  --0010011011001111    0010011011010000    0010011011010001    0010011011010010    0010011011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09935 - 09939

  --0010011011010100    0010011011010101    0010011011010110    0010011011010111    0010011011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09940 - 09944

  --0010011011011001    0010011011011010    0010011011011011    0010011011011100    0010011011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09945 - 09949

  --0010011011011110    0010011011011111    0010011011100000    0010011011100001    0010011011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09950 - 09954

  --0010011011100011    0010011011100100    0010011011100101    0010011011100110    0010011011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09955 - 09959

  --0010011011101000    0010011011101001    0010011011101010    0010011011101011    0010011011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09960 - 09964

  --0010011011101101    0010011011101110    0010011011101111    0010011011110000    0010011011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09965 - 09969

  --0010011011110010    0010011011110011    0010011011110100    0010011011110101    0010011011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09970 - 09974

  --0010011011110111    0010011011111000    0010011011111001    0010011011111010    0010011011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09975 - 09979

  --0010011011111100    0010011011111101    0010011011111110    0010011011111111    0010011100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09980 - 09984

  --0010011100000001    0010011100000010    0010011100000011    0010011100000100    0010011100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09985 - 09989

  --0010011100000110    0010011100000111    0010011100001000    0010011100001001    0010011100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09990 - 09994

  --0010011100001011    0010011100001100    0010011100001101    0010011100001110    0010011100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 09995 - 09999

  --0010011100010000    0010011100010001    0010011100010010    0010011100010011    0010011100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10000 - 10004

  --0010011100010101    0010011100010110    0010011100010111    0010011100011000    0010011100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10005 - 10009

  --0010011100011010    0010011100011011    0010011100011100    0010011100011101    0010011100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10010 - 10014

  --0010011100011111    0010011100100000    0010011100100001    0010011100100010    0010011100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10015 - 10019

  --0010011100100100    0010011100100101    0010011100100110    0010011100100111    0010011100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10020 - 10024

  --0010011100101001    0010011100101010    0010011100101011    0010011100101100    0010011100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10025 - 10029

  --0010011100101110    0010011100101111    0010011100110000    0010011100110001    0010011100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10030 - 10034

  --0010011100110011    0010011100110100    0010011100110101    0010011100110110    0010011100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10035 - 10039

  --0010011100111000    0010011100111001    0010011100111010    0010011100111011    0010011100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10040 - 10044

  --0010011100111101    0010011100111110    0010011100111111    0010011101000000    0010011101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10045 - 10049

  --0010011101000010    0010011101000011    0010011101000100    0010011101000101    0010011101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10050 - 10054

  --0010011101000111    0010011101001000    0010011101001001    0010011101001010    0010011101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10055 - 10059

  --0010011101001100    0010011101001101    0010011101001110    0010011101001111    0010011101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10060 - 10064

  --0010011101010001    0010011101010010    0010011101010011    0010011101010100    0010011101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10065 - 10069

  --0010011101010110    0010011101010111    0010011101011000    0010011101011001    0010011101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10070 - 10074

  --0010011101011011    0010011101011100    0010011101011101    0010011101011110    0010011101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10075 - 10079

  --0010011101100000    0010011101100001    0010011101100010    0010011101100011    0010011101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10080 - 10084

  --0010011101100101    0010011101100110    0010011101100111    0010011101101000    0010011101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10085 - 10089

  --0010011101101010    0010011101101011    0010011101101100    0010011101101101    0010011101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10090 - 10094

  --0010011101101111    0010011101110000    0010011101110001    0010011101110010    0010011101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10095 - 10099

  --0010011101110100    0010011101110101    0010011101110110    0010011101110111    0010011101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10100 - 10104

  --0010011101111001    0010011101111010    0010011101111011    0010011101111100    0010011101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10105 - 10109

  --0010011101111110    0010011101111111    0010011110000000    0010011110000001    0010011110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10110 - 10114

  --0010011110000011    0010011110000100    0010011110000101    0010011110000110    0010011110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10115 - 10119

  --0010011110001000    0010011110001001    0010011110001010    0010011110001011    0010011110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10120 - 10124

  --0010011110001101    0010011110001110    0010011110001111    0010011110010000    0010011110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10125 - 10129

  --0010011110010010    0010011110010011    0010011110010100    0010011110010101    0010011110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10130 - 10134

  --0010011110010111    0010011110011000    0010011110011001    0010011110011010    0010011110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10135 - 10139

  --0010011110011100    0010011110011101    0010011110011110    0010011110011111    0010011110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10140 - 10144

  --0010011110100001    0010011110100010    0010011110100011    0010011110100100    0010011110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10145 - 10149

  --0010011110100110    0010011110100111    0010011110101000    0010011110101001    0010011110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10150 - 10154

  --0010011110101011    0010011110101100    0010011110101101    0010011110101110    0010011110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10155 - 10159

  --0010011110110000    0010011110110001    0010011110110010    0010011110110011    0010011110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10160 - 10164

  --0010011110110101    0010011110110110    0010011110110111    0010011110111000    0010011110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10165 - 10169

  --0010011110111010    0010011110111011    0010011110111100    0010011110111101    0010011110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10170 - 10174

  --0010011110111111    0010011111000000    0010011111000001    0010011111000010    0010011111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10175 - 10179

  --0010011111000100    0010011111000101    0010011111000110    0010011111000111    0010011111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10180 - 10184

  --0010011111001001    0010011111001010    0010011111001011    0010011111001100    0010011111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10185 - 10189

  --0010011111001110    0010011111001111    0010011111010000    0010011111010001    0010011111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10190 - 10194

  --0010011111010011    0010011111010100    0010011111010101    0010011111010110    0010011111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10195 - 10199

  --0010011111011000    0010011111011001    0010011111011010    0010011111011011    0010011111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10200 - 10204

  --0010011111011101    0010011111011110    0010011111011111    0010011111100000    0010011111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10205 - 10209

  --0010011111100010    0010011111100011    0010011111100100    0010011111100101    0010011111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10210 - 10214

  --0010011111100111    0010011111101000    0010011111101001    0010011111101010    0010011111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10215 - 10219

  --0010011111101100    0010011111101101    0010011111101110    0010011111101111    0010011111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10220 - 10224

  --0010011111110001    0010011111110010    0010011111110011    0010011111110100    0010011111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10225 - 10229

  --0010011111110110    0010011111110111    0010011111111000    0010011111111001    0010011111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10230 - 10234

  --0010011111111011    0010011111111100    0010011111111101    0010011111111110    0010011111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10235 - 10239

  --0010100000000000    0010100000000001    0010100000000010    0010100000000011    0010100000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10240 - 10244

  --0010100000000101    0010100000000110    0010100000000111    0010100000001000    0010100000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10245 - 10249

  --0010100000001010    0010100000001011    0010100000001100    0010100000001101    0010100000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10250 - 10254

  --0010100000001111    0010100000010000    0010100000010001    0010100000010010    0010100000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10255 - 10259

  --0010100000010100    0010100000010101    0010100000010110    0010100000010111    0010100000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10260 - 10264

  --0010100000011001    0010100000011010    0010100000011011    0010100000011100    0010100000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10265 - 10269

  --0010100000011110    0010100000011111    0010100000100000    0010100000100001    0010100000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10270 - 10274

  --0010100000100011    0010100000100100    0010100000100101    0010100000100110    0010100000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10275 - 10279

  --0010100000101000    0010100000101001    0010100000101010    0010100000101011    0010100000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10280 - 10284

  --0010100000101101    0010100000101110    0010100000101111    0010100000110000    0010100000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10285 - 10289

  --0010100000110010    0010100000110011    0010100000110100    0010100000110101    0010100000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10290 - 10294

  --0010100000110111    0010100000111000    0010100000111001    0010100000111010    0010100000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10295 - 10299

  --0010100000111100    0010100000111101    0010100000111110    0010100000111111    0010100001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10300 - 10304

  --0010100001000001    0010100001000010    0010100001000011    0010100001000100    0010100001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10305 - 10309

  --0010100001000110    0010100001000111    0010100001001000    0010100001001001    0010100001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10310 - 10314

  --0010100001001011    0010100001001100    0010100001001101    0010100001001110    0010100001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10315 - 10319

  --0010100001010000    0010100001010001    0010100001010010    0010100001010011    0010100001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10320 - 10324

  --0010100001010101    0010100001010110    0010100001010111    0010100001011000    0010100001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10325 - 10329

  --0010100001011010    0010100001011011    0010100001011100    0010100001011101    0010100001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10330 - 10334

  --0010100001011111    0010100001100000    0010100001100001    0010100001100010    0010100001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10335 - 10339

  --0010100001100100    0010100001100101    0010100001100110    0010100001100111    0010100001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10340 - 10344

  --0010100001101001    0010100001101010    0010100001101011    0010100001101100    0010100001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10345 - 10349

  --0010100001101110    0010100001101111    0010100001110000    0010100001110001    0010100001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10350 - 10354

  --0010100001110011    0010100001110100    0010100001110101    0010100001110110    0010100001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10355 - 10359

  --0010100001111000    0010100001111001    0010100001111010    0010100001111011    0010100001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10360 - 10364

  --0010100001111101    0010100001111110    0010100001111111    0010100010000000    0010100010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10365 - 10369

  --0010100010000010    0010100010000011    0010100010000100    0010100010000101    0010100010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10370 - 10374

  --0010100010000111    0010100010001000    0010100010001001    0010100010001010    0010100010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10375 - 10379

  --0010100010001100    0010100010001101    0010100010001110    0010100010001111    0010100010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10380 - 10384

  --0010100010010001    0010100010010010    0010100010010011    0010100010010100    0010100010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10385 - 10389

  --0010100010010110    0010100010010111    0010100010011000    0010100010011001    0010100010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10390 - 10394

  --0010100010011011    0010100010011100    0010100010011101    0010100010011110    0010100010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10395 - 10399

  --0010100010100000    0010100010100001    0010100010100010    0010100010100011    0010100010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10400 - 10404

  --0010100010100101    0010100010100110    0010100010100111    0010100010101000    0010100010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10405 - 10409

  --0010100010101010    0010100010101011    0010100010101100    0010100010101101    0010100010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10410 - 10414

  --0010100010101111    0010100010110000    0010100010110001    0010100010110010    0010100010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10415 - 10419

  --0010100010110100    0010100010110101    0010100010110110    0010100010110111    0010100010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10420 - 10424

  --0010100010111001    0010100010111010    0010100010111011    0010100010111100    0010100010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10425 - 10429

  --0010100010111110    0010100010111111    0010100011000000    0010100011000001    0010100011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10430 - 10434

  --0010100011000011    0010100011000100    0010100011000101    0010100011000110    0010100011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10435 - 10439

  --0010100011001000    0010100011001001    0010100011001010    0010100011001011    0010100011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10440 - 10444

  --0010100011001101    0010100011001110    0010100011001111    0010100011010000    0010100011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10445 - 10449

  --0010100011010010    0010100011010011    0010100011010100    0010100011010101    0010100011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10450 - 10454

  --0010100011010111    0010100011011000    0010100011011001    0010100011011010    0010100011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10455 - 10459

  --0010100011011100    0010100011011101    0010100011011110    0010100011011111    0010100011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10460 - 10464

  --0010100011100001    0010100011100010    0010100011100011    0010100011100100    0010100011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10465 - 10469

  --0010100011100110    0010100011100111    0010100011101000    0010100011101001    0010100011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10470 - 10474

  --0010100011101011    0010100011101100    0010100011101101    0010100011101110    0010100011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10475 - 10479

  --0010100011110000    0010100011110001    0010100011110010    0010100011110011    0010100011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10480 - 10484

  --0010100011110101    0010100011110110    0010100011110111    0010100011111000    0010100011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10485 - 10489

  --0010100011111010    0010100011111011    0010100011111100    0010100011111101    0010100011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10490 - 10494

  --0010100011111111    0010100100000000    0010100100000001    0010100100000010    0010100100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10495 - 10499

  --0010100100000100    0010100100000101    0010100100000110    0010100100000111    0010100100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10500 - 10504

  --0010100100001001    0010100100001010    0010100100001011    0010100100001100    0010100100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10505 - 10509

  --0010100100001110    0010100100001111    0010100100010000    0010100100010001    0010100100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10510 - 10514

  --0010100100010011    0010100100010100    0010100100010101    0010100100010110    0010100100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10515 - 10519

  --0010100100011000    0010100100011001    0010100100011010    0010100100011011    0010100100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10520 - 10524

  --0010100100011101    0010100100011110    0010100100011111    0010100100100000    0010100100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10525 - 10529

  --0010100100100010    0010100100100011    0010100100100100    0010100100100101    0010100100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10530 - 10534

  --0010100100100111    0010100100101000    0010100100101001    0010100100101010    0010100100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10535 - 10539

  --0010100100101100    0010100100101101    0010100100101110    0010100100101111    0010100100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10540 - 10544

  --0010100100110001    0010100100110010    0010100100110011    0010100100110100    0010100100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10545 - 10549

  --0010100100110110    0010100100110111    0010100100111000    0010100100111001    0010100100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10550 - 10554

  --0010100100111011    0010100100111100    0010100100111101    0010100100111110    0010100100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10555 - 10559

  --0010100101000000    0010100101000001    0010100101000010    0010100101000011    0010100101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10560 - 10564

  --0010100101000101    0010100101000110    0010100101000111    0010100101001000    0010100101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10565 - 10569

  --0010100101001010    0010100101001011    0010100101001100    0010100101001101    0010100101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10570 - 10574

  --0010100101001111    0010100101010000    0010100101010001    0010100101010010    0010100101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10575 - 10579

  --0010100101010100    0010100101010101    0010100101010110    0010100101010111    0010100101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10580 - 10584

  --0010100101011001    0010100101011010    0010100101011011    0010100101011100    0010100101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10585 - 10589

  --0010100101011110    0010100101011111    0010100101100000    0010100101100001    0010100101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10590 - 10594

  --0010100101100011    0010100101100100    0010100101100101    0010100101100110    0010100101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10595 - 10599

  --0010100101101000    0010100101101001    0010100101101010    0010100101101011    0010100101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10600 - 10604

  --0010100101101101    0010100101101110    0010100101101111    0010100101110000    0010100101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10605 - 10609

  --0010100101110010    0010100101110011    0010100101110100    0010100101110101    0010100101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10610 - 10614

  --0010100101110111    0010100101111000    0010100101111001    0010100101111010    0010100101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10615 - 10619

  --0010100101111100    0010100101111101    0010100101111110    0010100101111111    0010100110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10620 - 10624

  --0010100110000001    0010100110000010    0010100110000011    0010100110000100    0010100110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10625 - 10629

  --0010100110000110    0010100110000111    0010100110001000    0010100110001001    0010100110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10630 - 10634

  --0010100110001011    0010100110001100    0010100110001101    0010100110001110    0010100110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10635 - 10639

  --0010100110010000    0010100110010001    0010100110010010    0010100110010011    0010100110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10640 - 10644

  --0010100110010101    0010100110010110    0010100110010111    0010100110011000    0010100110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10645 - 10649

  --0010100110011010    0010100110011011    0010100110011100    0010100110011101    0010100110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10650 - 10654

  --0010100110011111    0010100110100000    0010100110100001    0010100110100010    0010100110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10655 - 10659

  --0010100110100100    0010100110100101    0010100110100110    0010100110100111    0010100110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10660 - 10664

  --0010100110101001    0010100110101010    0010100110101011    0010100110101100    0010100110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10665 - 10669

  --0010100110101110    0010100110101111    0010100110110000    0010100110110001    0010100110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10670 - 10674

  --0010100110110011    0010100110110100    0010100110110101    0010100110110110    0010100110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10675 - 10679

  --0010100110111000    0010100110111001    0010100110111010    0010100110111011    0010100110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10680 - 10684

  --0010100110111101    0010100110111110    0010100110111111    0010100111000000    0010100111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10685 - 10689

  --0010100111000010    0010100111000011    0010100111000100    0010100111000101    0010100111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10690 - 10694

  --0010100111000111    0010100111001000    0010100111001001    0010100111001010    0010100111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10695 - 10699

  --0010100111001100    0010100111001101    0010100111001110    0010100111001111    0010100111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10700 - 10704

  --0010100111010001    0010100111010010    0010100111010011    0010100111010100    0010100111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10705 - 10709

  --0010100111010110    0010100111010111    0010100111011000    0010100111011001    0010100111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10710 - 10714

  --0010100111011011    0010100111011100    0010100111011101    0010100111011110    0010100111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10715 - 10719

  --0010100111100000    0010100111100001    0010100111100010    0010100111100011    0010100111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10720 - 10724

  --0010100111100101    0010100111100110    0010100111100111    0010100111101000    0010100111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10725 - 10729

  --0010100111101010    0010100111101011    0010100111101100    0010100111101101    0010100111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10730 - 10734

  --0010100111101111    0010100111110000    0010100111110001    0010100111110010    0010100111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10735 - 10739

  --0010100111110100    0010100111110101    0010100111110110    0010100111110111    0010100111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10740 - 10744

  --0010100111111001    0010100111111010    0010100111111011    0010100111111100    0010100111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10745 - 10749

  --0010100111111110    0010100111111111    0010101000000000    0010101000000001    0010101000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10750 - 10754

  --0010101000000011    0010101000000100    0010101000000101    0010101000000110    0010101000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10755 - 10759

  --0010101000001000    0010101000001001    0010101000001010    0010101000001011    0010101000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10760 - 10764

  --0010101000001101    0010101000001110    0010101000001111    0010101000010000    0010101000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10765 - 10769

  --0010101000010010    0010101000010011    0010101000010100    0010101000010101    0010101000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10770 - 10774

  --0010101000010111    0010101000011000    0010101000011001    0010101000011010    0010101000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10775 - 10779

  --0010101000011100    0010101000011101    0010101000011110    0010101000011111    0010101000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10780 - 10784

  --0010101000100001    0010101000100010    0010101000100011    0010101000100100    0010101000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10785 - 10789

  --0010101000100110    0010101000100111    0010101000101000    0010101000101001    0010101000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10790 - 10794

  --0010101000101011    0010101000101100    0010101000101101    0010101000101110    0010101000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10795 - 10799

  --0010101000110000    0010101000110001    0010101000110010    0010101000110011    0010101000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10800 - 10804

  --0010101000110101    0010101000110110    0010101000110111    0010101000111000    0010101000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10805 - 10809

  --0010101000111010    0010101000111011    0010101000111100    0010101000111101    0010101000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10810 - 10814

  --0010101000111111    0010101001000000    0010101001000001    0010101001000010    0010101001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10815 - 10819

  --0010101001000100    0010101001000101    0010101001000110    0010101001000111    0010101001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10820 - 10824

  --0010101001001001    0010101001001010    0010101001001011    0010101001001100    0010101001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10825 - 10829

  --0010101001001110    0010101001001111    0010101001010000    0010101001010001    0010101001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10830 - 10834

  --0010101001010011    0010101001010100    0010101001010101    0010101001010110    0010101001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10835 - 10839

  --0010101001011000    0010101001011001    0010101001011010    0010101001011011    0010101001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10840 - 10844

  --0010101001011101    0010101001011110    0010101001011111    0010101001100000    0010101001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10845 - 10849

  --0010101001100010    0010101001100011    0010101001100100    0010101001100101    0010101001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10850 - 10854

  --0010101001100111    0010101001101000    0010101001101001    0010101001101010    0010101001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10855 - 10859

  --0010101001101100    0010101001101101    0010101001101110    0010101001101111    0010101001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10860 - 10864

  --0010101001110001    0010101001110010    0010101001110011    0010101001110100    0010101001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10865 - 10869

  --0010101001110110    0010101001110111    0010101001111000    0010101001111001    0010101001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10870 - 10874

  --0010101001111011    0010101001111100    0010101001111101    0010101001111110    0010101001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10875 - 10879

  --0010101010000000    0010101010000001    0010101010000010    0010101010000011    0010101010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10880 - 10884

  --0010101010000101    0010101010000110    0010101010000111    0010101010001000    0010101010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10885 - 10889

  --0010101010001010    0010101010001011    0010101010001100    0010101010001101    0010101010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10890 - 10894

  --0010101010001111    0010101010010000    0010101010010001    0010101010010010    0010101010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10895 - 10899

  --0010101010010100    0010101010010101    0010101010010110    0010101010010111    0010101010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10900 - 10904

  --0010101010011001    0010101010011010    0010101010011011    0010101010011100    0010101010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10905 - 10909

  --0010101010011110    0010101010011111    0010101010100000    0010101010100001    0010101010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10910 - 10914

  --0010101010100011    0010101010100100    0010101010100101    0010101010100110    0010101010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10915 - 10919

  --0010101010101000    0010101010101001    0010101010101010    0010101010101011    0010101010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10920 - 10924

  --0010101010101101    0010101010101110    0010101010101111    0010101010110000    0010101010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10925 - 10929

  --0010101010110010    0010101010110011    0010101010110100    0010101010110101    0010101010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10930 - 10934

  --0010101010110111    0010101010111000    0010101010111001    0010101010111010    0010101010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10935 - 10939

  --0010101010111100    0010101010111101    0010101010111110    0010101010111111    0010101011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10940 - 10944

  --0010101011000001    0010101011000010    0010101011000011    0010101011000100    0010101011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10945 - 10949

  --0010101011000110    0010101011000111    0010101011001000    0010101011001001    0010101011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10950 - 10954

  --0010101011001011    0010101011001100    0010101011001101    0010101011001110    0010101011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10955 - 10959

  --0010101011010000    0010101011010001    0010101011010010    0010101011010011    0010101011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10960 - 10964

  --0010101011010101    0010101011010110    0010101011010111    0010101011011000    0010101011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10965 - 10969

  --0010101011011010    0010101011011011    0010101011011100    0010101011011101    0010101011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10970 - 10974

  --0010101011011111    0010101011100000    0010101011100001    0010101011100010    0010101011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10975 - 10979

  --0010101011100100    0010101011100101    0010101011100110    0010101011100111    0010101011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10980 - 10984

  --0010101011101001    0010101011101010    0010101011101011    0010101011101100    0010101011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10985 - 10989

  --0010101011101110    0010101011101111    0010101011110000    0010101011110001    0010101011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10990 - 10994

  --0010101011110011    0010101011110100    0010101011110101    0010101011110110    0010101011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 10995 - 10999

  --0010101011111000    0010101011111001    0010101011111010    0010101011111011    0010101011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11000 - 11004

  --0010101011111101    0010101011111110    0010101011111111    0010101100000000    0010101100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11005 - 11009

  --0010101100000010    0010101100000011    0010101100000100    0010101100000101    0010101100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11010 - 11014

  --0010101100000111    0010101100001000    0010101100001001    0010101100001010    0010101100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11015 - 11019

  --0010101100001100    0010101100001101    0010101100001110    0010101100001111    0010101100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11020 - 11024

  --0010101100010001    0010101100010010    0010101100010011    0010101100010100    0010101100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11025 - 11029

  --0010101100010110    0010101100010111    0010101100011000    0010101100011001    0010101100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11030 - 11034

  --0010101100011011    0010101100011100    0010101100011101    0010101100011110    0010101100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11035 - 11039

  --0010101100100000    0010101100100001    0010101100100010    0010101100100011    0010101100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11040 - 11044

  --0010101100100101    0010101100100110    0010101100100111    0010101100101000    0010101100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11045 - 11049

  --0010101100101010    0010101100101011    0010101100101100    0010101100101101    0010101100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11050 - 11054

  --0010101100101111    0010101100110000    0010101100110001    0010101100110010    0010101100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11055 - 11059

  --0010101100110100    0010101100110101    0010101100110110    0010101100110111    0010101100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11060 - 11064

  --0010101100111001    0010101100111010    0010101100111011    0010101100111100    0010101100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11065 - 11069

  --0010101100111110    0010101100111111    0010101101000000    0010101101000001    0010101101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11070 - 11074

  --0010101101000011    0010101101000100    0010101101000101    0010101101000110    0010101101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11075 - 11079

  --0010101101001000    0010101101001001    0010101101001010    0010101101001011    0010101101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11080 - 11084

  --0010101101001101    0010101101001110    0010101101001111    0010101101010000    0010101101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11085 - 11089

  --0010101101010010    0010101101010011    0010101101010100    0010101101010101    0010101101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11090 - 11094

  --0010101101010111    0010101101011000    0010101101011001    0010101101011010    0010101101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11095 - 11099

  --0010101101011100    0010101101011101    0010101101011110    0010101101011111    0010101101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11100 - 11104

  --0010101101100001    0010101101100010    0010101101100011    0010101101100100    0010101101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11105 - 11109

  --0010101101100110    0010101101100111    0010101101101000    0010101101101001    0010101101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11110 - 11114

  --0010101101101011    0010101101101100    0010101101101101    0010101101101110    0010101101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11115 - 11119

  --0010101101110000    0010101101110001    0010101101110010    0010101101110011    0010101101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11120 - 11124

  --0010101101110101    0010101101110110    0010101101110111    0010101101111000    0010101101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11125 - 11129

  --0010101101111010    0010101101111011    0010101101111100    0010101101111101    0010101101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11130 - 11134

  --0010101101111111    0010101110000000    0010101110000001    0010101110000010    0010101110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11135 - 11139

  --0010101110000100    0010101110000101    0010101110000110    0010101110000111    0010101110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11140 - 11144

  --0010101110001001    0010101110001010    0010101110001011    0010101110001100    0010101110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11145 - 11149

  --0010101110001110    0010101110001111    0010101110010000    0010101110010001    0010101110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11150 - 11154

  --0010101110010011    0010101110010100    0010101110010101    0010101110010110    0010101110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11155 - 11159

  --0010101110011000    0010101110011001    0010101110011010    0010101110011011    0010101110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11160 - 11164

  --0010101110011101    0010101110011110    0010101110011111    0010101110100000    0010101110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11165 - 11169

  --0010101110100010    0010101110100011    0010101110100100    0010101110100101    0010101110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11170 - 11174

  --0010101110100111    0010101110101000    0010101110101001    0010101110101010    0010101110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11175 - 11179

  --0010101110101100    0010101110101101    0010101110101110    0010101110101111    0010101110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11180 - 11184

  --0010101110110001    0010101110110010    0010101110110011    0010101110110100    0010101110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11185 - 11189

  --0010101110110110    0010101110110111    0010101110111000    0010101110111001    0010101110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11190 - 11194

  --0010101110111011    0010101110111100    0010101110111101    0010101110111110    0010101110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11195 - 11199

  --0010101111000000    0010101111000001    0010101111000010    0010101111000011    0010101111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11200 - 11204

  --0010101111000101    0010101111000110    0010101111000111    0010101111001000    0010101111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11205 - 11209

  --0010101111001010    0010101111001011    0010101111001100    0010101111001101    0010101111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11210 - 11214

  --0010101111001111    0010101111010000    0010101111010001    0010101111010010    0010101111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11215 - 11219

  --0010101111010100    0010101111010101    0010101111010110    0010101111010111    0010101111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11220 - 11224

  --0010101111011001    0010101111011010    0010101111011011    0010101111011100    0010101111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11225 - 11229

  --0010101111011110    0010101111011111    0010101111100000    0010101111100001    0010101111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11230 - 11234

  --0010101111100011    0010101111100100    0010101111100101    0010101111100110    0010101111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11235 - 11239

  --0010101111101000    0010101111101001    0010101111101010    0010101111101011    0010101111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11240 - 11244

  --0010101111101101    0010101111101110    0010101111101111    0010101111110000    0010101111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11245 - 11249

  --0010101111110010    0010101111110011    0010101111110100    0010101111110101    0010101111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11250 - 11254

  --0010101111110111    0010101111111000    0010101111111001    0010101111111010    0010101111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11255 - 11259

  --0010101111111100    0010101111111101    0010101111111110    0010101111111111    0010110000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11260 - 11264

  --0010110000000001    0010110000000010    0010110000000011    0010110000000100    0010110000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11265 - 11269

  --0010110000000110    0010110000000111    0010110000001000    0010110000001001    0010110000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11270 - 11274

  --0010110000001011    0010110000001100    0010110000001101    0010110000001110    0010110000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11275 - 11279

  --0010110000010000    0010110000010001    0010110000010010    0010110000010011    0010110000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11280 - 11284

  --0010110000010101    0010110000010110    0010110000010111    0010110000011000    0010110000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11285 - 11289

  --0010110000011010    0010110000011011    0010110000011100    0010110000011101    0010110000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11290 - 11294

  --0010110000011111    0010110000100000    0010110000100001    0010110000100010    0010110000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11295 - 11299

  --0010110000100100    0010110000100101    0010110000100110    0010110000100111    0010110000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11300 - 11304

  --0010110000101001    0010110000101010    0010110000101011    0010110000101100    0010110000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11305 - 11309

  --0010110000101110    0010110000101111    0010110000110000    0010110000110001    0010110000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11310 - 11314

  --0010110000110011    0010110000110100    0010110000110101    0010110000110110    0010110000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11315 - 11319

  --0010110000111000    0010110000111001    0010110000111010    0010110000111011    0010110000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11320 - 11324

  --0010110000111101    0010110000111110    0010110000111111    0010110001000000    0010110001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11325 - 11329

  --0010110001000010    0010110001000011    0010110001000100    0010110001000101    0010110001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11330 - 11334

  --0010110001000111    0010110001001000    0010110001001001    0010110001001010    0010110001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11335 - 11339

  --0010110001001100    0010110001001101    0010110001001110    0010110001001111    0010110001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11340 - 11344

  --0010110001010001    0010110001010010    0010110001010011    0010110001010100    0010110001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11345 - 11349

  --0010110001010110    0010110001010111    0010110001011000    0010110001011001    0010110001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11350 - 11354

  --0010110001011011    0010110001011100    0010110001011101    0010110001011110    0010110001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11355 - 11359

  --0010110001100000    0010110001100001    0010110001100010    0010110001100011    0010110001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11360 - 11364

  --0010110001100101    0010110001100110    0010110001100111    0010110001101000    0010110001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11365 - 11369

  --0010110001101010    0010110001101011    0010110001101100    0010110001101101    0010110001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11370 - 11374

  --0010110001101111    0010110001110000    0010110001110001    0010110001110010    0010110001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11375 - 11379

  --0010110001110100    0010110001110101    0010110001110110    0010110001110111    0010110001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11380 - 11384

  --0010110001111001    0010110001111010    0010110001111011    0010110001111100    0010110001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11385 - 11389

  --0010110001111110    0010110001111111    0010110010000000    0010110010000001    0010110010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11390 - 11394

  --0010110010000011    0010110010000100    0010110010000101    0010110010000110    0010110010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11395 - 11399

  --0010110010001000    0010110010001001    0010110010001010    0010110010001011    0010110010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11400 - 11404

  --0010110010001101    0010110010001110    0010110010001111    0010110010010000    0010110010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11405 - 11409

  --0010110010010010    0010110010010011    0010110010010100    0010110010010101    0010110010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11410 - 11414

  --0010110010010111    0010110010011000    0010110010011001    0010110010011010    0010110010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11415 - 11419

  --0010110010011100    0010110010011101    0010110010011110    0010110010011111    0010110010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11420 - 11424

  --0010110010100001    0010110010100010    0010110010100011    0010110010100100    0010110010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11425 - 11429

  --0010110010100110    0010110010100111    0010110010101000    0010110010101001    0010110010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11430 - 11434

  --0010110010101011    0010110010101100    0010110010101101    0010110010101110    0010110010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11435 - 11439

  --0010110010110000    0010110010110001    0010110010110010    0010110010110011    0010110010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11440 - 11444

  --0010110010110101    0010110010110110    0010110010110111    0010110010111000    0010110010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11445 - 11449

  --0010110010111010    0010110010111011    0010110010111100    0010110010111101    0010110010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11450 - 11454

  --0010110010111111    0010110011000000    0010110011000001    0010110011000010    0010110011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11455 - 11459

  --0010110011000100    0010110011000101    0010110011000110    0010110011000111    0010110011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11460 - 11464

  --0010110011001001    0010110011001010    0010110011001011    0010110011001100    0010110011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11465 - 11469

  --0010110011001110    0010110011001111    0010110011010000    0010110011010001    0010110011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11470 - 11474

  --0010110011010011    0010110011010100    0010110011010101    0010110011010110    0010110011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11475 - 11479

  --0010110011011000    0010110011011001    0010110011011010    0010110011011011    0010110011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11480 - 11484

  --0010110011011101    0010110011011110    0010110011011111    0010110011100000    0010110011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11485 - 11489

  --0010110011100010    0010110011100011    0010110011100100    0010110011100101    0010110011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11490 - 11494

  --0010110011100111    0010110011101000    0010110011101001    0010110011101010    0010110011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11495 - 11499

  --0010110011101100    0010110011101101    0010110011101110    0010110011101111    0010110011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11500 - 11504

  --0010110011110001    0010110011110010    0010110011110011    0010110011110100    0010110011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11505 - 11509

  --0010110011110110    0010110011110111    0010110011111000    0010110011111001    0010110011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11510 - 11514

  --0010110011111011    0010110011111100    0010110011111101    0010110011111110    0010110011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11515 - 11519

  --0010110100000000    0010110100000001    0010110100000010    0010110100000011    0010110100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11520 - 11524

  --0010110100000101    0010110100000110    0010110100000111    0010110100001000    0010110100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11525 - 11529

  --0010110100001010    0010110100001011    0010110100001100    0010110100001101    0010110100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11530 - 11534

  --0010110100001111    0010110100010000    0010110100010001    0010110100010010    0010110100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11535 - 11539

  --0010110100010100    0010110100010101    0010110100010110    0010110100010111    0010110100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11540 - 11544

  --0010110100011001    0010110100011010    0010110100011011    0010110100011100    0010110100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11545 - 11549

  --0010110100011110    0010110100011111    0010110100100000    0010110100100001    0010110100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11550 - 11554

  --0010110100100011    0010110100100100    0010110100100101    0010110100100110    0010110100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11555 - 11559

  --0010110100101000    0010110100101001    0010110100101010    0010110100101011    0010110100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11560 - 11564

  --0010110100101101    0010110100101110    0010110100101111    0010110100110000    0010110100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11565 - 11569

  --0010110100110010    0010110100110011    0010110100110100    0010110100110101    0010110100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11570 - 11574

  --0010110100110111    0010110100111000    0010110100111001    0010110100111010    0010110100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11575 - 11579

  --0010110100111100    0010110100111101    0010110100111110    0010110100111111    0010110101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11580 - 11584

  --0010110101000001    0010110101000010    0010110101000011    0010110101000100    0010110101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11585 - 11589

  --0010110101000110    0010110101000111    0010110101001000    0010110101001001    0010110101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11590 - 11594

  --0010110101001011    0010110101001100    0010110101001101    0010110101001110    0010110101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11595 - 11599

  --0010110101010000    0010110101010001    0010110101010010    0010110101010011    0010110101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11600 - 11604

  --0010110101010101    0010110101010110    0010110101010111    0010110101011000    0010110101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11605 - 11609

  --0010110101011010    0010110101011011    0010110101011100    0010110101011101    0010110101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11610 - 11614

  --0010110101011111    0010110101100000    0010110101100001    0010110101100010    0010110101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11615 - 11619

  --0010110101100100    0010110101100101    0010110101100110    0010110101100111    0010110101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11620 - 11624

  --0010110101101001    0010110101101010    0010110101101011    0010110101101100    0010110101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11625 - 11629

  --0010110101101110    0010110101101111    0010110101110000    0010110101110001    0010110101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11630 - 11634

  --0010110101110011    0010110101110100    0010110101110101    0010110101110110    0010110101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11635 - 11639

  --0010110101111000    0010110101111001    0010110101111010    0010110101111011    0010110101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11640 - 11644

  --0010110101111101    0010110101111110    0010110101111111    0010110110000000    0010110110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11645 - 11649

  --0010110110000010    0010110110000011    0010110110000100    0010110110000101    0010110110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11650 - 11654

  --0010110110000111    0010110110001000    0010110110001001    0010110110001010    0010110110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11655 - 11659

  --0010110110001100    0010110110001101    0010110110001110    0010110110001111    0010110110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11660 - 11664

  --0010110110010001    0010110110010010    0010110110010011    0010110110010100    0010110110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11665 - 11669

  --0010110110010110    0010110110010111    0010110110011000    0010110110011001    0010110110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11670 - 11674

  --0010110110011011    0010110110011100    0010110110011101    0010110110011110    0010110110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11675 - 11679

  --0010110110100000    0010110110100001    0010110110100010    0010110110100011    0010110110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11680 - 11684

  --0010110110100101    0010110110100110    0010110110100111    0010110110101000    0010110110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11685 - 11689

  --0010110110101010    0010110110101011    0010110110101100    0010110110101101    0010110110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11690 - 11694

  --0010110110101111    0010110110110000    0010110110110001    0010110110110010    0010110110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11695 - 11699

  --0010110110110100    0010110110110101    0010110110110110    0010110110110111    0010110110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11700 - 11704

  --0010110110111001    0010110110111010    0010110110111011    0010110110111100    0010110110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11705 - 11709

  --0010110110111110    0010110110111111    0010110111000000    0010110111000001    0010110111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11710 - 11714

  --0010110111000011    0010110111000100    0010110111000101    0010110111000110    0010110111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11715 - 11719

  --0010110111001000    0010110111001001    0010110111001010    0010110111001011    0010110111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11720 - 11724

  --0010110111001101    0010110111001110    0010110111001111    0010110111010000    0010110111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11725 - 11729

  --0010110111010010    0010110111010011    0010110111010100    0010110111010101    0010110111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11730 - 11734

  --0010110111010111    0010110111011000    0010110111011001    0010110111011010    0010110111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11735 - 11739

  --0010110111011100    0010110111011101    0010110111011110    0010110111011111    0010110111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11740 - 11744

  --0010110111100001    0010110111100010    0010110111100011    0010110111100100    0010110111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11745 - 11749

  --0010110111100110    0010110111100111    0010110111101000    0010110111101001    0010110111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11750 - 11754

  --0010110111101011    0010110111101100    0010110111101101    0010110111101110    0010110111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11755 - 11759

  --0010110111110000    0010110111110001    0010110111110010    0010110111110011    0010110111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11760 - 11764

  --0010110111110101    0010110111110110    0010110111110111    0010110111111000    0010110111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11765 - 11769

  --0010110111111010    0010110111111011    0010110111111100    0010110111111101    0010110111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11770 - 11774

  --0010110111111111    0010111000000000    0010111000000001    0010111000000010    0010111000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11775 - 11779

  --0010111000000100    0010111000000101    0010111000000110    0010111000000111    0010111000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11780 - 11784

  --0010111000001001    0010111000001010    0010111000001011    0010111000001100    0010111000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11785 - 11789

  --0010111000001110    0010111000001111    0010111000010000    0010111000010001    0010111000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11790 - 11794

  --0010111000010011    0010111000010100    0010111000010101    0010111000010110    0010111000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11795 - 11799

  --0010111000011000    0010111000011001    0010111000011010    0010111000011011    0010111000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11800 - 11804

  --0010111000011101    0010111000011110    0010111000011111    0010111000100000    0010111000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11805 - 11809

  --0010111000100010    0010111000100011    0010111000100100    0010111000100101    0010111000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11810 - 11814

  --0010111000100111    0010111000101000    0010111000101001    0010111000101010    0010111000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11815 - 11819

  --0010111000101100    0010111000101101    0010111000101110    0010111000101111    0010111000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11820 - 11824

  --0010111000110001    0010111000110010    0010111000110011    0010111000110100    0010111000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11825 - 11829

  --0010111000110110    0010111000110111    0010111000111000    0010111000111001    0010111000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11830 - 11834

  --0010111000111011    0010111000111100    0010111000111101    0010111000111110    0010111000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11835 - 11839

  --0010111001000000    0010111001000001    0010111001000010    0010111001000011    0010111001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11840 - 11844

  --0010111001000101    0010111001000110    0010111001000111    0010111001001000    0010111001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11845 - 11849

  --0010111001001010    0010111001001011    0010111001001100    0010111001001101    0010111001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11850 - 11854

  --0010111001001111    0010111001010000    0010111001010001    0010111001010010    0010111001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11855 - 11859

  --0010111001010100    0010111001010101    0010111001010110    0010111001010111    0010111001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11860 - 11864

  --0010111001011001    0010111001011010    0010111001011011    0010111001011100    0010111001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11865 - 11869

  --0010111001011110    0010111001011111    0010111001100000    0010111001100001    0010111001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11870 - 11874

  --0010111001100011    0010111001100100    0010111001100101    0010111001100110    0010111001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11875 - 11879

  --0010111001101000    0010111001101001    0010111001101010    0010111001101011    0010111001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11880 - 11884

  --0010111001101101    0010111001101110    0010111001101111    0010111001110000    0010111001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11885 - 11889

  --0010111001110010    0010111001110011    0010111001110100    0010111001110101    0010111001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11890 - 11894

  --0010111001110111    0010111001111000    0010111001111001    0010111001111010    0010111001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11895 - 11899

  --0010111001111100    0010111001111101    0010111001111110    0010111001111111    0010111010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11900 - 11904

  --0010111010000001    0010111010000010    0010111010000011    0010111010000100    0010111010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11905 - 11909

  --0010111010000110    0010111010000111    0010111010001000    0010111010001001    0010111010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11910 - 11914

  --0010111010001011    0010111010001100    0010111010001101    0010111010001110    0010111010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11915 - 11919

  --0010111010010000    0010111010010001    0010111010010010    0010111010010011    0010111010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11920 - 11924

  --0010111010010101    0010111010010110    0010111010010111    0010111010011000    0010111010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11925 - 11929

  --0010111010011010    0010111010011011    0010111010011100    0010111010011101    0010111010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11930 - 11934

  --0010111010011111    0010111010100000    0010111010100001    0010111010100010    0010111010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11935 - 11939

  --0010111010100100    0010111010100101    0010111010100110    0010111010100111    0010111010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11940 - 11944

  --0010111010101001    0010111010101010    0010111010101011    0010111010101100    0010111010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11945 - 11949

  --0010111010101110    0010111010101111    0010111010110000    0010111010110001    0010111010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11950 - 11954

  --0010111010110011    0010111010110100    0010111010110101    0010111010110110    0010111010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11955 - 11959

  --0010111010111000    0010111010111001    0010111010111010    0010111010111011    0010111010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11960 - 11964

  --0010111010111101    0010111010111110    0010111010111111    0010111011000000    0010111011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11965 - 11969

  --0010111011000010    0010111011000011    0010111011000100    0010111011000101    0010111011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11970 - 11974

  --0010111011000111    0010111011001000    0010111011001001    0010111011001010    0010111011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11975 - 11979

  --0010111011001100    0010111011001101    0010111011001110    0010111011001111    0010111011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11980 - 11984

  --0010111011010001    0010111011010010    0010111011010011    0010111011010100    0010111011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11985 - 11989

  --0010111011010110    0010111011010111    0010111011011000    0010111011011001    0010111011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11990 - 11994

  --0010111011011011    0010111011011100    0010111011011101    0010111011011110    0010111011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 11995 - 11999

  --0010111011100000    0010111011100001    0010111011100010    0010111011100011    0010111011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12000 - 12004

  --0010111011100101    0010111011100110    0010111011100111    0010111011101000    0010111011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12005 - 12009

  --0010111011101010    0010111011101011    0010111011101100    0010111011101101    0010111011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12010 - 12014

  --0010111011101111    0010111011110000    0010111011110001    0010111011110010    0010111011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12015 - 12019

  --0010111011110100    0010111011110101    0010111011110110    0010111011110111    0010111011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12020 - 12024

  --0010111011111001    0010111011111010    0010111011111011    0010111011111100    0010111011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12025 - 12029

  --0010111011111110    0010111011111111    0010111100000000    0010111100000001    0010111100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12030 - 12034

  --0010111100000011    0010111100000100    0010111100000101    0010111100000110    0010111100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12035 - 12039

  --0010111100001000    0010111100001001    0010111100001010    0010111100001011    0010111100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12040 - 12044

  --0010111100001101    0010111100001110    0010111100001111    0010111100010000    0010111100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12045 - 12049

  --0010111100010010    0010111100010011    0010111100010100    0010111100010101    0010111100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12050 - 12054

  --0010111100010111    0010111100011000    0010111100011001    0010111100011010    0010111100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12055 - 12059

  --0010111100011100    0010111100011101    0010111100011110    0010111100011111    0010111100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12060 - 12064

  --0010111100100001    0010111100100010    0010111100100011    0010111100100100    0010111100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12065 - 12069

  --0010111100100110    0010111100100111    0010111100101000    0010111100101001    0010111100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12070 - 12074

  --0010111100101011    0010111100101100    0010111100101101    0010111100101110    0010111100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12075 - 12079

  --0010111100110000    0010111100110001    0010111100110010    0010111100110011    0010111100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12080 - 12084

  --0010111100110101    0010111100110110    0010111100110111    0010111100111000    0010111100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12085 - 12089

  --0010111100111010    0010111100111011    0010111100111100    0010111100111101    0010111100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12090 - 12094

  --0010111100111111    0010111101000000    0010111101000001    0010111101000010    0010111101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12095 - 12099

  --0010111101000100    0010111101000101    0010111101000110    0010111101000111    0010111101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12100 - 12104

  --0010111101001001    0010111101001010    0010111101001011    0010111101001100    0010111101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12105 - 12109

  --0010111101001110    0010111101001111    0010111101010000    0010111101010001    0010111101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12110 - 12114

  --0010111101010011    0010111101010100    0010111101010101    0010111101010110    0010111101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12115 - 12119

  --0010111101011000    0010111101011001    0010111101011010    0010111101011011    0010111101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12120 - 12124

  --0010111101011101    0010111101011110    0010111101011111    0010111101100000    0010111101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12125 - 12129

  --0010111101100010    0010111101100011    0010111101100100    0010111101100101    0010111101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12130 - 12134

  --0010111101100111    0010111101101000    0010111101101001    0010111101101010    0010111101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12135 - 12139

  --0010111101101100    0010111101101101    0010111101101110    0010111101101111    0010111101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12140 - 12144

  --0010111101110001    0010111101110010    0010111101110011    0010111101110100    0010111101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12145 - 12149

  --0010111101110110    0010111101110111    0010111101111000    0010111101111001    0010111101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12150 - 12154

  --0010111101111011    0010111101111100    0010111101111101    0010111101111110    0010111101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12155 - 12159

  --0010111110000000    0010111110000001    0010111110000010    0010111110000011    0010111110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12160 - 12164

  --0010111110000101    0010111110000110    0010111110000111    0010111110001000    0010111110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12165 - 12169

  --0010111110001010    0010111110001011    0010111110001100    0010111110001101    0010111110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12170 - 12174

  --0010111110001111    0010111110010000    0010111110010001    0010111110010010    0010111110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12175 - 12179

  --0010111110010100    0010111110010101    0010111110010110    0010111110010111    0010111110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12180 - 12184

  --0010111110011001    0010111110011010    0010111110011011    0010111110011100    0010111110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12185 - 12189

  --0010111110011110    0010111110011111    0010111110100000    0010111110100001    0010111110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12190 - 12194

  --0010111110100011    0010111110100100    0010111110100101    0010111110100110    0010111110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12195 - 12199

  --0010111110101000    0010111110101001    0010111110101010    0010111110101011    0010111110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12200 - 12204

  --0010111110101101    0010111110101110    0010111110101111    0010111110110000    0010111110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12205 - 12209

  --0010111110110010    0010111110110011    0010111110110100    0010111110110101    0010111110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12210 - 12214

  --0010111110110111    0010111110111000    0010111110111001    0010111110111010    0010111110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12215 - 12219

  --0010111110111100    0010111110111101    0010111110111110    0010111110111111    0010111111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12220 - 12224

  --0010111111000001    0010111111000010    0010111111000011    0010111111000100    0010111111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12225 - 12229

  --0010111111000110    0010111111000111    0010111111001000    0010111111001001    0010111111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12230 - 12234

  --0010111111001011    0010111111001100    0010111111001101    0010111111001110    0010111111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12235 - 12239

  --0010111111010000    0010111111010001    0010111111010010    0010111111010011    0010111111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12240 - 12244

  --0010111111010101    0010111111010110    0010111111010111    0010111111011000    0010111111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12245 - 12249

  --0010111111011010    0010111111011011    0010111111011100    0010111111011101    0010111111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12250 - 12254

  --0010111111011111    0010111111100000    0010111111100001    0010111111100010    0010111111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12255 - 12259

  --0010111111100100    0010111111100101    0010111111100110    0010111111100111    0010111111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12260 - 12264

  --0010111111101001    0010111111101010    0010111111101011    0010111111101100    0010111111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12265 - 12269

  --0010111111101110    0010111111101111    0010111111110000    0010111111110001    0010111111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12270 - 12274

  --0010111111110011    0010111111110100    0010111111110101    0010111111110110    0010111111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12275 - 12279

  --0010111111111000    0010111111111001    0010111111111010    0010111111111011    0010111111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12280 - 12284

  --0010111111111101    0010111111111110    0010111111111111    0011000000000000    0011000000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12285 - 12289

  --0011000000000010    0011000000000011    0011000000000100    0011000000000101    0011000000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12290 - 12294

  --0011000000000111    0011000000001000    0011000000001001    0011000000001010    0011000000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12295 - 12299

  --0011000000001100    0011000000001101    0011000000001110    0011000000001111    0011000000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12300 - 12304

  --0011000000010001    0011000000010010    0011000000010011    0011000000010100    0011000000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12305 - 12309

  --0011000000010110    0011000000010111    0011000000011000    0011000000011001    0011000000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12310 - 12314

  --0011000000011011    0011000000011100    0011000000011101    0011000000011110    0011000000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12315 - 12319

  --0011000000100000    0011000000100001    0011000000100010    0011000000100011    0011000000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12320 - 12324

  --0011000000100101    0011000000100110    0011000000100111    0011000000101000    0011000000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12325 - 12329

  --0011000000101010    0011000000101011    0011000000101100    0011000000101101    0011000000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12330 - 12334

  --0011000000101111    0011000000110000    0011000000110001    0011000000110010    0011000000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12335 - 12339

  --0011000000110100    0011000000110101    0011000000110110    0011000000110111    0011000000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12340 - 12344

  --0011000000111001    0011000000111010    0011000000111011    0011000000111100    0011000000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12345 - 12349

  --0011000000111110    0011000000111111    0011000001000000    0011000001000001    0011000001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12350 - 12354

  --0011000001000011    0011000001000100    0011000001000101    0011000001000110    0011000001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12355 - 12359

  --0011000001001000    0011000001001001    0011000001001010    0011000001001011    0011000001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12360 - 12364

  --0011000001001101    0011000001001110    0011000001001111    0011000001010000    0011000001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12365 - 12369

  --0011000001010010    0011000001010011    0011000001010100    0011000001010101    0011000001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12370 - 12374

  --0011000001010111    0011000001011000    0011000001011001    0011000001011010    0011000001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12375 - 12379

  --0011000001011100    0011000001011101    0011000001011110    0011000001011111    0011000001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12380 - 12384

  --0011000001100001    0011000001100010    0011000001100011    0011000001100100    0011000001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12385 - 12389

  --0011000001100110    0011000001100111    0011000001101000    0011000001101001    0011000001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12390 - 12394

  --0011000001101011    0011000001101100    0011000001101101    0011000001101110    0011000001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12395 - 12399

  --0011000001110000    0011000001110001    0011000001110010    0011000001110011    0011000001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12400 - 12404

  --0011000001110101    0011000001110110    0011000001110111    0011000001111000    0011000001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12405 - 12409

  --0011000001111010    0011000001111011    0011000001111100    0011000001111101    0011000001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12410 - 12414

  --0011000001111111    0011000010000000    0011000010000001    0011000010000010    0011000010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12415 - 12419

  --0011000010000100    0011000010000101    0011000010000110    0011000010000111    0011000010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12420 - 12424

  --0011000010001001    0011000010001010    0011000010001011    0011000010001100    0011000010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12425 - 12429

  --0011000010001110    0011000010001111    0011000010010000    0011000010010001    0011000010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12430 - 12434

  --0011000010010011    0011000010010100    0011000010010101    0011000010010110    0011000010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12435 - 12439

  --0011000010011000    0011000010011001    0011000010011010    0011000010011011    0011000010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12440 - 12444

  --0011000010011101    0011000010011110    0011000010011111    0011000010100000    0011000010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12445 - 12449

  --0011000010100010    0011000010100011    0011000010100100    0011000010100101    0011000010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12450 - 12454

  --0011000010100111    0011000010101000    0011000010101001    0011000010101010    0011000010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12455 - 12459

  --0011000010101100    0011000010101101    0011000010101110    0011000010101111    0011000010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12460 - 12464

  --0011000010110001    0011000010110010    0011000010110011    0011000010110100    0011000010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12465 - 12469

  --0011000010110110    0011000010110111    0011000010111000    0011000010111001    0011000010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12470 - 12474

  --0011000010111011    0011000010111100    0011000010111101    0011000010111110    0011000010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12475 - 12479

  --0011000011000000    0011000011000001    0011000011000010    0011000011000011    0011000011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12480 - 12484

  --0011000011000101    0011000011000110    0011000011000111    0011000011001000    0011000011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12485 - 12489

  --0011000011001010    0011000011001011    0011000011001100    0011000011001101    0011000011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12490 - 12494

  --0011000011001111    0011000011010000    0011000011010001    0011000011010010    0011000011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12495 - 12499

  --0011000011010100    0011000011010101    0011000011010110    0011000011010111    0011000011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12500 - 12504

  --0011000011011001    0011000011011010    0011000011011011    0011000011011100    0011000011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12505 - 12509

  --0011000011011110    0011000011011111    0011000011100000    0011000011100001    0011000011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12510 - 12514

  --0011000011100011    0011000011100100    0011000011100101    0011000011100110    0011000011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12515 - 12519

  --0011000011101000    0011000011101001    0011000011101010    0011000011101011    0011000011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12520 - 12524

  --0011000011101101    0011000011101110    0011000011101111    0011000011110000    0011000011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12525 - 12529

  --0011000011110010    0011000011110011    0011000011110100    0011000011110101    0011000011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12530 - 12534

  --0011000011110111    0011000011111000    0011000011111001    0011000011111010    0011000011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12535 - 12539

  --0011000011111100    0011000011111101    0011000011111110    0011000011111111    0011000100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12540 - 12544

  --0011000100000001    0011000100000010    0011000100000011    0011000100000100    0011000100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12545 - 12549

  --0011000100000110    0011000100000111    0011000100001000    0011000100001001    0011000100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12550 - 12554

  --0011000100001011    0011000100001100    0011000100001101    0011000100001110    0011000100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12555 - 12559

  --0011000100010000    0011000100010001    0011000100010010    0011000100010011    0011000100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12560 - 12564

  --0011000100010101    0011000100010110    0011000100010111    0011000100011000    0011000100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12565 - 12569

  --0011000100011010    0011000100011011    0011000100011100    0011000100011101    0011000100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12570 - 12574

  --0011000100011111    0011000100100000    0011000100100001    0011000100100010    0011000100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12575 - 12579

  --0011000100100100    0011000100100101    0011000100100110    0011000100100111    0011000100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12580 - 12584

  --0011000100101001    0011000100101010    0011000100101011    0011000100101100    0011000100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12585 - 12589

  --0011000100101110    0011000100101111    0011000100110000    0011000100110001    0011000100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12590 - 12594

  --0011000100110011    0011000100110100    0011000100110101    0011000100110110    0011000100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12595 - 12599

  --0011000100111000    0011000100111001    0011000100111010    0011000100111011    0011000100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12600 - 12604

  --0011000100111101    0011000100111110    0011000100111111    0011000101000000    0011000101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12605 - 12609

  --0011000101000010    0011000101000011    0011000101000100    0011000101000101    0011000101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12610 - 12614

  --0011000101000111    0011000101001000    0011000101001001    0011000101001010    0011000101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12615 - 12619

  --0011000101001100    0011000101001101    0011000101001110    0011000101001111    0011000101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12620 - 12624

  --0011000101010001    0011000101010010    0011000101010011    0011000101010100    0011000101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12625 - 12629

  --0011000101010110    0011000101010111    0011000101011000    0011000101011001    0011000101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12630 - 12634

  --0011000101011011    0011000101011100    0011000101011101    0011000101011110    0011000101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12635 - 12639

  --0011000101100000    0011000101100001    0011000101100010    0011000101100011    0011000101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12640 - 12644

  --0011000101100101    0011000101100110    0011000101100111    0011000101101000    0011000101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12645 - 12649

  --0011000101101010    0011000101101011    0011000101101100    0011000101101101    0011000101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12650 - 12654

  --0011000101101111    0011000101110000    0011000101110001    0011000101110010    0011000101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12655 - 12659

  --0011000101110100    0011000101110101    0011000101110110    0011000101110111    0011000101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12660 - 12664

  --0011000101111001    0011000101111010    0011000101111011    0011000101111100    0011000101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12665 - 12669

  --0011000101111110    0011000101111111    0011000110000000    0011000110000001    0011000110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12670 - 12674

  --0011000110000011    0011000110000100    0011000110000101    0011000110000110    0011000110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12675 - 12679

  --0011000110001000    0011000110001001    0011000110001010    0011000110001011    0011000110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12680 - 12684

  --0011000110001101    0011000110001110    0011000110001111    0011000110010000    0011000110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12685 - 12689

  --0011000110010010    0011000110010011    0011000110010100    0011000110010101    0011000110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12690 - 12694

  --0011000110010111    0011000110011000    0011000110011001    0011000110011010    0011000110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12695 - 12699

  --0011000110011100    0011000110011101    0011000110011110    0011000110011111    0011000110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12700 - 12704

  --0011000110100001    0011000110100010    0011000110100011    0011000110100100    0011000110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12705 - 12709

  --0011000110100110    0011000110100111    0011000110101000    0011000110101001    0011000110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12710 - 12714

  --0011000110101011    0011000110101100    0011000110101101    0011000110101110    0011000110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12715 - 12719

  --0011000110110000    0011000110110001    0011000110110010    0011000110110011    0011000110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12720 - 12724

  --0011000110110101    0011000110110110    0011000110110111    0011000110111000    0011000110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12725 - 12729

  --0011000110111010    0011000110111011    0011000110111100    0011000110111101    0011000110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12730 - 12734

  --0011000110111111    0011000111000000    0011000111000001    0011000111000010    0011000111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12735 - 12739

  --0011000111000100    0011000111000101    0011000111000110    0011000111000111    0011000111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12740 - 12744

  --0011000111001001    0011000111001010    0011000111001011    0011000111001100    0011000111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12745 - 12749

  --0011000111001110    0011000111001111    0011000111010000    0011000111010001    0011000111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12750 - 12754

  --0011000111010011    0011000111010100    0011000111010101    0011000111010110    0011000111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12755 - 12759

  --0011000111011000    0011000111011001    0011000111011010    0011000111011011    0011000111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12760 - 12764

  --0011000111011101    0011000111011110    0011000111011111    0011000111100000    0011000111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12765 - 12769

  --0011000111100010    0011000111100011    0011000111100100    0011000111100101    0011000111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12770 - 12774

  --0011000111100111    0011000111101000    0011000111101001    0011000111101010    0011000111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12775 - 12779

  --0011000111101100    0011000111101101    0011000111101110    0011000111101111    0011000111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12780 - 12784

  --0011000111110001    0011000111110010    0011000111110011    0011000111110100    0011000111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12785 - 12789

  --0011000111110110    0011000111110111    0011000111111000    0011000111111001    0011000111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12790 - 12794

  --0011000111111011    0011000111111100    0011000111111101    0011000111111110    0011000111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12795 - 12799

  --0011001000000000    0011001000000001    0011001000000010    0011001000000011    0011001000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12800 - 12804

  --0011001000000101    0011001000000110    0011001000000111    0011001000001000    0011001000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12805 - 12809

  --0011001000001010    0011001000001011    0011001000001100    0011001000001101    0011001000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12810 - 12814

  --0011001000001111    0011001000010000    0011001000010001    0011001000010010    0011001000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12815 - 12819

  --0011001000010100    0011001000010101    0011001000010110    0011001000010111    0011001000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12820 - 12824

  --0011001000011001    0011001000011010    0011001000011011    0011001000011100    0011001000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12825 - 12829

  --0011001000011110    0011001000011111    0011001000100000    0011001000100001    0011001000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12830 - 12834

  --0011001000100011    0011001000100100    0011001000100101    0011001000100110    0011001000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12835 - 12839

  --0011001000101000    0011001000101001    0011001000101010    0011001000101011    0011001000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12840 - 12844

  --0011001000101101    0011001000101110    0011001000101111    0011001000110000    0011001000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12845 - 12849

  --0011001000110010    0011001000110011    0011001000110100    0011001000110101    0011001000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12850 - 12854

  --0011001000110111    0011001000111000    0011001000111001    0011001000111010    0011001000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12855 - 12859

  --0011001000111100    0011001000111101    0011001000111110    0011001000111111    0011001001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12860 - 12864

  --0011001001000001    0011001001000010    0011001001000011    0011001001000100    0011001001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12865 - 12869

  --0011001001000110    0011001001000111    0011001001001000    0011001001001001    0011001001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12870 - 12874

  --0011001001001011    0011001001001100    0011001001001101    0011001001001110    0011001001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12875 - 12879

  --0011001001010000    0011001001010001    0011001001010010    0011001001010011    0011001001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12880 - 12884

  --0011001001010101    0011001001010110    0011001001010111    0011001001011000    0011001001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12885 - 12889

  --0011001001011010    0011001001011011    0011001001011100    0011001001011101    0011001001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12890 - 12894

  --0011001001011111    0011001001100000    0011001001100001    0011001001100010    0011001001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12895 - 12899

  --0011001001100100    0011001001100101    0011001001100110    0011001001100111    0011001001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12900 - 12904

  --0011001001101001    0011001001101010    0011001001101011    0011001001101100    0011001001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12905 - 12909

  --0011001001101110    0011001001101111    0011001001110000    0011001001110001    0011001001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12910 - 12914

  --0011001001110011    0011001001110100    0011001001110101    0011001001110110    0011001001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12915 - 12919

  --0011001001111000    0011001001111001    0011001001111010    0011001001111011    0011001001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12920 - 12924

  --0011001001111101    0011001001111110    0011001001111111    0011001010000000    0011001010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12925 - 12929

  --0011001010000010    0011001010000011    0011001010000100    0011001010000101    0011001010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12930 - 12934

  --0011001010000111    0011001010001000    0011001010001001    0011001010001010    0011001010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12935 - 12939

  --0011001010001100    0011001010001101    0011001010001110    0011001010001111    0011001010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12940 - 12944

  --0011001010010001    0011001010010010    0011001010010011    0011001010010100    0011001010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12945 - 12949

  --0011001010010110    0011001010010111    0011001010011000    0011001010011001    0011001010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12950 - 12954

  --0011001010011011    0011001010011100    0011001010011101    0011001010011110    0011001010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12955 - 12959

  --0011001010100000    0011001010100001    0011001010100010    0011001010100011    0011001010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12960 - 12964

  --0011001010100101    0011001010100110    0011001010100111    0011001010101000    0011001010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12965 - 12969

  --0011001010101010    0011001010101011    0011001010101100    0011001010101101    0011001010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12970 - 12974

  --0011001010101111    0011001010110000    0011001010110001    0011001010110010    0011001010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12975 - 12979

  --0011001010110100    0011001010110101    0011001010110110    0011001010110111    0011001010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12980 - 12984

  --0011001010111001    0011001010111010    0011001010111011    0011001010111100    0011001010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12985 - 12989

  --0011001010111110    0011001010111111    0011001011000000    0011001011000001    0011001011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12990 - 12994

  --0011001011000011    0011001011000100    0011001011000101    0011001011000110    0011001011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 12995 - 12999

  --0011001011001000    0011001011001001    0011001011001010    0011001011001011    0011001011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13000 - 13004

  --0011001011001101    0011001011001110    0011001011001111    0011001011010000    0011001011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13005 - 13009

  --0011001011010010    0011001011010011    0011001011010100    0011001011010101    0011001011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13010 - 13014

  --0011001011010111    0011001011011000    0011001011011001    0011001011011010    0011001011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13015 - 13019

  --0011001011011100    0011001011011101    0011001011011110    0011001011011111    0011001011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13020 - 13024

  --0011001011100001    0011001011100010    0011001011100011    0011001011100100    0011001011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13025 - 13029

  --0011001011100110    0011001011100111    0011001011101000    0011001011101001    0011001011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13030 - 13034

  --0011001011101011    0011001011101100    0011001011101101    0011001011101110    0011001011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13035 - 13039

  --0011001011110000    0011001011110001    0011001011110010    0011001011110011    0011001011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13040 - 13044

  --0011001011110101    0011001011110110    0011001011110111    0011001011111000    0011001011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13045 - 13049

  --0011001011111010    0011001011111011    0011001011111100    0011001011111101    0011001011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13050 - 13054

  --0011001011111111    0011001100000000    0011001100000001    0011001100000010    0011001100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13055 - 13059

  --0011001100000100    0011001100000101    0011001100000110    0011001100000111    0011001100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13060 - 13064

  --0011001100001001    0011001100001010    0011001100001011    0011001100001100    0011001100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13065 - 13069

  --0011001100001110    0011001100001111    0011001100010000    0011001100010001    0011001100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13070 - 13074

  --0011001100010011    0011001100010100    0011001100010101    0011001100010110    0011001100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13075 - 13079

  --0011001100011000    0011001100011001    0011001100011010    0011001100011011    0011001100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13080 - 13084

  --0011001100011101    0011001100011110    0011001100011111    0011001100100000    0011001100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13085 - 13089

  --0011001100100010    0011001100100011    0011001100100100    0011001100100101    0011001100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13090 - 13094

  --0011001100100111    0011001100101000    0011001100101001    0011001100101010    0011001100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13095 - 13099

  --0011001100101100    0011001100101101    0011001100101110    0011001100101111    0011001100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13100 - 13104

  --0011001100110001    0011001100110010    0011001100110011    0011001100110100    0011001100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13105 - 13109

  --0011001100110110    0011001100110111    0011001100111000    0011001100111001    0011001100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13110 - 13114

  --0011001100111011    0011001100111100    0011001100111101    0011001100111110    0011001100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13115 - 13119

  --0011001101000000    0011001101000001    0011001101000010    0011001101000011    0011001101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13120 - 13124

  --0011001101000101    0011001101000110    0011001101000111    0011001101001000    0011001101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13125 - 13129

  --0011001101001010    0011001101001011    0011001101001100    0011001101001101    0011001101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13130 - 13134

  --0011001101001111    0011001101010000    0011001101010001    0011001101010010    0011001101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13135 - 13139

  --0011001101010100    0011001101010101    0011001101010110    0011001101010111    0011001101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13140 - 13144

  --0011001101011001    0011001101011010    0011001101011011    0011001101011100    0011001101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13145 - 13149

  --0011001101011110    0011001101011111    0011001101100000    0011001101100001    0011001101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13150 - 13154

  --0011001101100011    0011001101100100    0011001101100101    0011001101100110    0011001101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13155 - 13159

  --0011001101101000    0011001101101001    0011001101101010    0011001101101011    0011001101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13160 - 13164

  --0011001101101101    0011001101101110    0011001101101111    0011001101110000    0011001101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13165 - 13169

  --0011001101110010    0011001101110011    0011001101110100    0011001101110101    0011001101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13170 - 13174

  --0011001101110111    0011001101111000    0011001101111001    0011001101111010    0011001101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13175 - 13179

  --0011001101111100    0011001101111101    0011001101111110    0011001101111111    0011001110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13180 - 13184

  --0011001110000001    0011001110000010    0011001110000011    0011001110000100    0011001110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13185 - 13189

  --0011001110000110    0011001110000111    0011001110001000    0011001110001001    0011001110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13190 - 13194

  --0011001110001011    0011001110001100    0011001110001101    0011001110001110    0011001110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13195 - 13199

  --0011001110010000    0011001110010001    0011001110010010    0011001110010011    0011001110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13200 - 13204

  --0011001110010101    0011001110010110    0011001110010111    0011001110011000    0011001110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13205 - 13209

  --0011001110011010    0011001110011011    0011001110011100    0011001110011101    0011001110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13210 - 13214

  --0011001110011111    0011001110100000    0011001110100001    0011001110100010    0011001110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13215 - 13219

  --0011001110100100    0011001110100101    0011001110100110    0011001110100111    0011001110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13220 - 13224

  --0011001110101001    0011001110101010    0011001110101011    0011001110101100    0011001110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13225 - 13229

  --0011001110101110    0011001110101111    0011001110110000    0011001110110001    0011001110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13230 - 13234

  --0011001110110011    0011001110110100    0011001110110101    0011001110110110    0011001110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13235 - 13239

  --0011001110111000    0011001110111001    0011001110111010    0011001110111011    0011001110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13240 - 13244

  --0011001110111101    0011001110111110    0011001110111111    0011001111000000    0011001111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13245 - 13249

  --0011001111000010    0011001111000011    0011001111000100    0011001111000101    0011001111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13250 - 13254

  --0011001111000111    0011001111001000    0011001111001001    0011001111001010    0011001111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13255 - 13259

  --0011001111001100    0011001111001101    0011001111001110    0011001111001111    0011001111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13260 - 13264

  --0011001111010001    0011001111010010    0011001111010011    0011001111010100    0011001111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13265 - 13269

  --0011001111010110    0011001111010111    0011001111011000    0011001111011001    0011001111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13270 - 13274

  --0011001111011011    0011001111011100    0011001111011101    0011001111011110    0011001111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13275 - 13279

  --0011001111100000    0011001111100001    0011001111100010    0011001111100011    0011001111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13280 - 13284

  --0011001111100101    0011001111100110    0011001111100111    0011001111101000    0011001111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13285 - 13289

  --0011001111101010    0011001111101011    0011001111101100    0011001111101101    0011001111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13290 - 13294

  --0011001111101111    0011001111110000    0011001111110001    0011001111110010    0011001111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13295 - 13299

  --0011001111110100    0011001111110101    0011001111110110    0011001111110111    0011001111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13300 - 13304

  --0011001111111001    0011001111111010    0011001111111011    0011001111111100    0011001111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13305 - 13309

  --0011001111111110    0011001111111111    0011010000000000    0011010000000001    0011010000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13310 - 13314

  --0011010000000011    0011010000000100    0011010000000101    0011010000000110    0011010000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13315 - 13319

  --0011010000001000    0011010000001001    0011010000001010    0011010000001011    0011010000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13320 - 13324

  --0011010000001101    0011010000001110    0011010000001111    0011010000010000    0011010000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13325 - 13329

  --0011010000010010    0011010000010011    0011010000010100    0011010000010101    0011010000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13330 - 13334

  --0011010000010111    0011010000011000    0011010000011001    0011010000011010    0011010000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13335 - 13339

  --0011010000011100    0011010000011101    0011010000011110    0011010000011111    0011010000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13340 - 13344

  --0011010000100001    0011010000100010    0011010000100011    0011010000100100    0011010000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13345 - 13349

  --0011010000100110    0011010000100111    0011010000101000    0011010000101001    0011010000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13350 - 13354

  --0011010000101011    0011010000101100    0011010000101101    0011010000101110    0011010000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13355 - 13359

  --0011010000110000    0011010000110001    0011010000110010    0011010000110011    0011010000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13360 - 13364

  --0011010000110101    0011010000110110    0011010000110111    0011010000111000    0011010000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13365 - 13369

  --0011010000111010    0011010000111011    0011010000111100    0011010000111101    0011010000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13370 - 13374

  --0011010000111111    0011010001000000    0011010001000001    0011010001000010    0011010001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13375 - 13379

  --0011010001000100    0011010001000101    0011010001000110    0011010001000111    0011010001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13380 - 13384

  --0011010001001001    0011010001001010    0011010001001011    0011010001001100    0011010001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13385 - 13389

  --0011010001001110    0011010001001111    0011010001010000    0011010001010001    0011010001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13390 - 13394

  --0011010001010011    0011010001010100    0011010001010101    0011010001010110    0011010001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13395 - 13399

  --0011010001011000    0011010001011001    0011010001011010    0011010001011011    0011010001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13400 - 13404

  --0011010001011101    0011010001011110    0011010001011111    0011010001100000    0011010001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13405 - 13409

  --0011010001100010    0011010001100011    0011010001100100    0011010001100101    0011010001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13410 - 13414

  --0011010001100111    0011010001101000    0011010001101001    0011010001101010    0011010001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13415 - 13419

  --0011010001101100    0011010001101101    0011010001101110    0011010001101111    0011010001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13420 - 13424

  --0011010001110001    0011010001110010    0011010001110011    0011010001110100    0011010001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13425 - 13429

  --0011010001110110    0011010001110111    0011010001111000    0011010001111001    0011010001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13430 - 13434

  --0011010001111011    0011010001111100    0011010001111101    0011010001111110    0011010001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13435 - 13439

  --0011010010000000    0011010010000001    0011010010000010    0011010010000011    0011010010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13440 - 13444

  --0011010010000101    0011010010000110    0011010010000111    0011010010001000    0011010010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13445 - 13449

  --0011010010001010    0011010010001011    0011010010001100    0011010010001101    0011010010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13450 - 13454

  --0011010010001111    0011010010010000    0011010010010001    0011010010010010    0011010010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13455 - 13459

  --0011010010010100    0011010010010101    0011010010010110    0011010010010111    0011010010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13460 - 13464

  --0011010010011001    0011010010011010    0011010010011011    0011010010011100    0011010010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13465 - 13469

  --0011010010011110    0011010010011111    0011010010100000    0011010010100001    0011010010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13470 - 13474

  --0011010010100011    0011010010100100    0011010010100101    0011010010100110    0011010010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13475 - 13479

  --0011010010101000    0011010010101001    0011010010101010    0011010010101011    0011010010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13480 - 13484

  --0011010010101101    0011010010101110    0011010010101111    0011010010110000    0011010010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13485 - 13489

  --0011010010110010    0011010010110011    0011010010110100    0011010010110101    0011010010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13490 - 13494

  --0011010010110111    0011010010111000    0011010010111001    0011010010111010    0011010010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13495 - 13499

  --0011010010111100    0011010010111101    0011010010111110    0011010010111111    0011010011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13500 - 13504

  --0011010011000001    0011010011000010    0011010011000011    0011010011000100    0011010011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13505 - 13509

  --0011010011000110    0011010011000111    0011010011001000    0011010011001001    0011010011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13510 - 13514

  --0011010011001011    0011010011001100    0011010011001101    0011010011001110    0011010011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13515 - 13519

  --0011010011010000    0011010011010001    0011010011010010    0011010011010011    0011010011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13520 - 13524

  --0011010011010101    0011010011010110    0011010011010111    0011010011011000    0011010011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13525 - 13529

  --0011010011011010    0011010011011011    0011010011011100    0011010011011101    0011010011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13530 - 13534

  --0011010011011111    0011010011100000    0011010011100001    0011010011100010    0011010011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13535 - 13539

  --0011010011100100    0011010011100101    0011010011100110    0011010011100111    0011010011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13540 - 13544

  --0011010011101001    0011010011101010    0011010011101011    0011010011101100    0011010011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13545 - 13549

  --0011010011101110    0011010011101111    0011010011110000    0011010011110001    0011010011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13550 - 13554

  --0011010011110011    0011010011110100    0011010011110101    0011010011110110    0011010011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13555 - 13559

  --0011010011111000    0011010011111001    0011010011111010    0011010011111011    0011010011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13560 - 13564

  --0011010011111101    0011010011111110    0011010011111111    0011010100000000    0011010100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13565 - 13569

  --0011010100000010    0011010100000011    0011010100000100    0011010100000101    0011010100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13570 - 13574

  --0011010100000111    0011010100001000    0011010100001001    0011010100001010    0011010100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13575 - 13579

  --0011010100001100    0011010100001101    0011010100001110    0011010100001111    0011010100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13580 - 13584

  --0011010100010001    0011010100010010    0011010100010011    0011010100010100    0011010100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13585 - 13589

  --0011010100010110    0011010100010111    0011010100011000    0011010100011001    0011010100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13590 - 13594

  --0011010100011011    0011010100011100    0011010100011101    0011010100011110    0011010100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13595 - 13599

  --0011010100100000    0011010100100001    0011010100100010    0011010100100011    0011010100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13600 - 13604

  --0011010100100101    0011010100100110    0011010100100111    0011010100101000    0011010100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13605 - 13609

  --0011010100101010    0011010100101011    0011010100101100    0011010100101101    0011010100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13610 - 13614

  --0011010100101111    0011010100110000    0011010100110001    0011010100110010    0011010100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13615 - 13619

  --0011010100110100    0011010100110101    0011010100110110    0011010100110111    0011010100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13620 - 13624

  --0011010100111001    0011010100111010    0011010100111011    0011010100111100    0011010100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13625 - 13629

  --0011010100111110    0011010100111111    0011010101000000    0011010101000001    0011010101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13630 - 13634

  --0011010101000011    0011010101000100    0011010101000101    0011010101000110    0011010101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13635 - 13639

  --0011010101001000    0011010101001001    0011010101001010    0011010101001011    0011010101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13640 - 13644

  --0011010101001101    0011010101001110    0011010101001111    0011010101010000    0011010101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13645 - 13649

  --0011010101010010    0011010101010011    0011010101010100    0011010101010101    0011010101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13650 - 13654

  --0011010101010111    0011010101011000    0011010101011001    0011010101011010    0011010101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13655 - 13659

  --0011010101011100    0011010101011101    0011010101011110    0011010101011111    0011010101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13660 - 13664

  --0011010101100001    0011010101100010    0011010101100011    0011010101100100    0011010101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13665 - 13669

  --0011010101100110    0011010101100111    0011010101101000    0011010101101001    0011010101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13670 - 13674

  --0011010101101011    0011010101101100    0011010101101101    0011010101101110    0011010101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13675 - 13679

  --0011010101110000    0011010101110001    0011010101110010    0011010101110011    0011010101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13680 - 13684

  --0011010101110101    0011010101110110    0011010101110111    0011010101111000    0011010101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13685 - 13689

  --0011010101111010    0011010101111011    0011010101111100    0011010101111101    0011010101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13690 - 13694

  --0011010101111111    0011010110000000    0011010110000001    0011010110000010    0011010110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13695 - 13699

  --0011010110000100    0011010110000101    0011010110000110    0011010110000111    0011010110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13700 - 13704

  --0011010110001001    0011010110001010    0011010110001011    0011010110001100    0011010110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13705 - 13709

  --0011010110001110    0011010110001111    0011010110010000    0011010110010001    0011010110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13710 - 13714

  --0011010110010011    0011010110010100    0011010110010101    0011010110010110    0011010110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13715 - 13719

  --0011010110011000    0011010110011001    0011010110011010    0011010110011011    0011010110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13720 - 13724

  --0011010110011101    0011010110011110    0011010110011111    0011010110100000    0011010110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13725 - 13729

  --0011010110100010    0011010110100011    0011010110100100    0011010110100101    0011010110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13730 - 13734

  --0011010110100111    0011010110101000    0011010110101001    0011010110101010    0011010110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13735 - 13739

  --0011010110101100    0011010110101101    0011010110101110    0011010110101111    0011010110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13740 - 13744

  --0011010110110001    0011010110110010    0011010110110011    0011010110110100    0011010110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13745 - 13749

  --0011010110110110    0011010110110111    0011010110111000    0011010110111001    0011010110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13750 - 13754

  --0011010110111011    0011010110111100    0011010110111101    0011010110111110    0011010110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13755 - 13759

  --0011010111000000    0011010111000001    0011010111000010    0011010111000011    0011010111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13760 - 13764

  --0011010111000101    0011010111000110    0011010111000111    0011010111001000    0011010111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13765 - 13769

  --0011010111001010    0011010111001011    0011010111001100    0011010111001101    0011010111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13770 - 13774

  --0011010111001111    0011010111010000    0011010111010001    0011010111010010    0011010111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13775 - 13779

  --0011010111010100    0011010111010101    0011010111010110    0011010111010111    0011010111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13780 - 13784

  --0011010111011001    0011010111011010    0011010111011011    0011010111011100    0011010111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13785 - 13789

  --0011010111011110    0011010111011111    0011010111100000    0011010111100001    0011010111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13790 - 13794

  --0011010111100011    0011010111100100    0011010111100101    0011010111100110    0011010111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13795 - 13799

  --0011010111101000    0011010111101001    0011010111101010    0011010111101011    0011010111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13800 - 13804

  --0011010111101101    0011010111101110    0011010111101111    0011010111110000    0011010111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13805 - 13809

  --0011010111110010    0011010111110011    0011010111110100    0011010111110101    0011010111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13810 - 13814

  --0011010111110111    0011010111111000    0011010111111001    0011010111111010    0011010111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13815 - 13819

  --0011010111111100    0011010111111101    0011010111111110    0011010111111111    0011011000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13820 - 13824

  --0011011000000001    0011011000000010    0011011000000011    0011011000000100    0011011000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13825 - 13829

  --0011011000000110    0011011000000111    0011011000001000    0011011000001001    0011011000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13830 - 13834

  --0011011000001011    0011011000001100    0011011000001101    0011011000001110    0011011000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13835 - 13839

  --0011011000010000    0011011000010001    0011011000010010    0011011000010011    0011011000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13840 - 13844

  --0011011000010101    0011011000010110    0011011000010111    0011011000011000    0011011000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13845 - 13849

  --0011011000011010    0011011000011011    0011011000011100    0011011000011101    0011011000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13850 - 13854

  --0011011000011111    0011011000100000    0011011000100001    0011011000100010    0011011000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13855 - 13859

  --0011011000100100    0011011000100101    0011011000100110    0011011000100111    0011011000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13860 - 13864

  --0011011000101001    0011011000101010    0011011000101011    0011011000101100    0011011000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13865 - 13869

  --0011011000101110    0011011000101111    0011011000110000    0011011000110001    0011011000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13870 - 13874

  --0011011000110011    0011011000110100    0011011000110101    0011011000110110    0011011000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13875 - 13879

  --0011011000111000    0011011000111001    0011011000111010    0011011000111011    0011011000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13880 - 13884

  --0011011000111101    0011011000111110    0011011000111111    0011011001000000    0011011001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13885 - 13889

  --0011011001000010    0011011001000011    0011011001000100    0011011001000101    0011011001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13890 - 13894

  --0011011001000111    0011011001001000    0011011001001001    0011011001001010    0011011001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13895 - 13899

  --0011011001001100    0011011001001101    0011011001001110    0011011001001111    0011011001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13900 - 13904

  --0011011001010001    0011011001010010    0011011001010011    0011011001010100    0011011001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13905 - 13909

  --0011011001010110    0011011001010111    0011011001011000    0011011001011001    0011011001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13910 - 13914

  --0011011001011011    0011011001011100    0011011001011101    0011011001011110    0011011001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13915 - 13919

  --0011011001100000    0011011001100001    0011011001100010    0011011001100011    0011011001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13920 - 13924

  --0011011001100101    0011011001100110    0011011001100111    0011011001101000    0011011001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13925 - 13929

  --0011011001101010    0011011001101011    0011011001101100    0011011001101101    0011011001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13930 - 13934

  --0011011001101111    0011011001110000    0011011001110001    0011011001110010    0011011001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13935 - 13939

  --0011011001110100    0011011001110101    0011011001110110    0011011001110111    0011011001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13940 - 13944

  --0011011001111001    0011011001111010    0011011001111011    0011011001111100    0011011001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13945 - 13949

  --0011011001111110    0011011001111111    0011011010000000    0011011010000001    0011011010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13950 - 13954

  --0011011010000011    0011011010000100    0011011010000101    0011011010000110    0011011010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13955 - 13959

  --0011011010001000    0011011010001001    0011011010001010    0011011010001011    0011011010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13960 - 13964

  --0011011010001101    0011011010001110    0011011010001111    0011011010010000    0011011010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13965 - 13969

  --0011011010010010    0011011010010011    0011011010010100    0011011010010101    0011011010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13970 - 13974

  --0011011010010111    0011011010011000    0011011010011001    0011011010011010    0011011010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13975 - 13979

  --0011011010011100    0011011010011101    0011011010011110    0011011010011111    0011011010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13980 - 13984

  --0011011010100001    0011011010100010    0011011010100011    0011011010100100    0011011010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13985 - 13989

  --0011011010100110    0011011010100111    0011011010101000    0011011010101001    0011011010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13990 - 13994

  --0011011010101011    0011011010101100    0011011010101101    0011011010101110    0011011010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 13995 - 13999

  --0011011010110000    0011011010110001    0011011010110010    0011011010110011    0011011010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14000 - 14004

  --0011011010110101    0011011010110110    0011011010110111    0011011010111000    0011011010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14005 - 14009

  --0011011010111010    0011011010111011    0011011010111100    0011011010111101    0011011010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14010 - 14014

  --0011011010111111    0011011011000000    0011011011000001    0011011011000010    0011011011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14015 - 14019

  --0011011011000100    0011011011000101    0011011011000110    0011011011000111    0011011011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14020 - 14024

  --0011011011001001    0011011011001010    0011011011001011    0011011011001100    0011011011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14025 - 14029

  --0011011011001110    0011011011001111    0011011011010000    0011011011010001    0011011011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14030 - 14034

  --0011011011010011    0011011011010100    0011011011010101    0011011011010110    0011011011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14035 - 14039

  --0011011011011000    0011011011011001    0011011011011010    0011011011011011    0011011011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14040 - 14044

  --0011011011011101    0011011011011110    0011011011011111    0011011011100000    0011011011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14045 - 14049

  --0011011011100010    0011011011100011    0011011011100100    0011011011100101    0011011011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14050 - 14054

  --0011011011100111    0011011011101000    0011011011101001    0011011011101010    0011011011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14055 - 14059

  --0011011011101100    0011011011101101    0011011011101110    0011011011101111    0011011011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14060 - 14064

  --0011011011110001    0011011011110010    0011011011110011    0011011011110100    0011011011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14065 - 14069

  --0011011011110110    0011011011110111    0011011011111000    0011011011111001    0011011011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14070 - 14074

  --0011011011111011    0011011011111100    0011011011111101    0011011011111110    0011011011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14075 - 14079

  --0011011100000000    0011011100000001    0011011100000010    0011011100000011    0011011100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14080 - 14084

  --0011011100000101    0011011100000110    0011011100000111    0011011100001000    0011011100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14085 - 14089

  --0011011100001010    0011011100001011    0011011100001100    0011011100001101    0011011100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14090 - 14094

  --0011011100001111    0011011100010000    0011011100010001    0011011100010010    0011011100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14095 - 14099

  --0011011100010100    0011011100010101    0011011100010110    0011011100010111    0011011100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14100 - 14104

  --0011011100011001    0011011100011010    0011011100011011    0011011100011100    0011011100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14105 - 14109

  --0011011100011110    0011011100011111    0011011100100000    0011011100100001    0011011100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14110 - 14114

  --0011011100100011    0011011100100100    0011011100100101    0011011100100110    0011011100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14115 - 14119

  --0011011100101000    0011011100101001    0011011100101010    0011011100101011    0011011100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14120 - 14124

  --0011011100101101    0011011100101110    0011011100101111    0011011100110000    0011011100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14125 - 14129

  --0011011100110010    0011011100110011    0011011100110100    0011011100110101    0011011100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14130 - 14134

  --0011011100110111    0011011100111000    0011011100111001    0011011100111010    0011011100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14135 - 14139

  --0011011100111100    0011011100111101    0011011100111110    0011011100111111    0011011101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14140 - 14144

  --0011011101000001    0011011101000010    0011011101000011    0011011101000100    0011011101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14145 - 14149

  --0011011101000110    0011011101000111    0011011101001000    0011011101001001    0011011101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14150 - 14154

  --0011011101001011    0011011101001100    0011011101001101    0011011101001110    0011011101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14155 - 14159

  --0011011101010000    0011011101010001    0011011101010010    0011011101010011    0011011101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14160 - 14164

  --0011011101010101    0011011101010110    0011011101010111    0011011101011000    0011011101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14165 - 14169

  --0011011101011010    0011011101011011    0011011101011100    0011011101011101    0011011101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14170 - 14174

  --0011011101011111    0011011101100000    0011011101100001    0011011101100010    0011011101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14175 - 14179

  --0011011101100100    0011011101100101    0011011101100110    0011011101100111    0011011101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14180 - 14184

  --0011011101101001    0011011101101010    0011011101101011    0011011101101100    0011011101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14185 - 14189

  --0011011101101110    0011011101101111    0011011101110000    0011011101110001    0011011101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14190 - 14194

  --0011011101110011    0011011101110100    0011011101110101    0011011101110110    0011011101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14195 - 14199

  --0011011101111000    0011011101111001    0011011101111010    0011011101111011    0011011101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14200 - 14204

  --0011011101111101    0011011101111110    0011011101111111    0011011110000000    0011011110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14205 - 14209

  --0011011110000010    0011011110000011    0011011110000100    0011011110000101    0011011110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14210 - 14214

  --0011011110000111    0011011110001000    0011011110001001    0011011110001010    0011011110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14215 - 14219

  --0011011110001100    0011011110001101    0011011110001110    0011011110001111    0011011110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14220 - 14224

  --0011011110010001    0011011110010010    0011011110010011    0011011110010100    0011011110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14225 - 14229

  --0011011110010110    0011011110010111    0011011110011000    0011011110011001    0011011110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14230 - 14234

  --0011011110011011    0011011110011100    0011011110011101    0011011110011110    0011011110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14235 - 14239

  --0011011110100000    0011011110100001    0011011110100010    0011011110100011    0011011110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14240 - 14244

  --0011011110100101    0011011110100110    0011011110100111    0011011110101000    0011011110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14245 - 14249

  --0011011110101010    0011011110101011    0011011110101100    0011011110101101    0011011110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14250 - 14254

  --0011011110101111    0011011110110000    0011011110110001    0011011110110010    0011011110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14255 - 14259

  --0011011110110100    0011011110110101    0011011110110110    0011011110110111    0011011110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14260 - 14264

  --0011011110111001    0011011110111010    0011011110111011    0011011110111100    0011011110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14265 - 14269

  --0011011110111110    0011011110111111    0011011111000000    0011011111000001    0011011111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14270 - 14274

  --0011011111000011    0011011111000100    0011011111000101    0011011111000110    0011011111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14275 - 14279

  --0011011111001000    0011011111001001    0011011111001010    0011011111001011    0011011111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14280 - 14284

  --0011011111001101    0011011111001110    0011011111001111    0011011111010000    0011011111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14285 - 14289

  --0011011111010010    0011011111010011    0011011111010100    0011011111010101    0011011111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14290 - 14294

  --0011011111010111    0011011111011000    0011011111011001    0011011111011010    0011011111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14295 - 14299

  --0011011111011100    0011011111011101    0011011111011110    0011011111011111    0011011111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14300 - 14304

  --0011011111100001    0011011111100010    0011011111100011    0011011111100100    0011011111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14305 - 14309

  --0011011111100110    0011011111100111    0011011111101000    0011011111101001    0011011111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14310 - 14314

  --0011011111101011    0011011111101100    0011011111101101    0011011111101110    0011011111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14315 - 14319

  --0011011111110000    0011011111110001    0011011111110010    0011011111110011    0011011111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14320 - 14324

  --0011011111110101    0011011111110110    0011011111110111    0011011111111000    0011011111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14325 - 14329

  --0011011111111010    0011011111111011    0011011111111100    0011011111111101    0011011111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14330 - 14334

  --0011011111111111    0011100000000000    0011100000000001    0011100000000010    0011100000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14335 - 14339

  --0011100000000100    0011100000000101    0011100000000110    0011100000000111    0011100000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14340 - 14344

  --0011100000001001    0011100000001010    0011100000001011    0011100000001100    0011100000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14345 - 14349

  --0011100000001110    0011100000001111    0011100000010000    0011100000010001    0011100000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14350 - 14354

  --0011100000010011    0011100000010100    0011100000010101    0011100000010110    0011100000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14355 - 14359

  --0011100000011000    0011100000011001    0011100000011010    0011100000011011    0011100000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14360 - 14364

  --0011100000011101    0011100000011110    0011100000011111    0011100000100000    0011100000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14365 - 14369

  --0011100000100010    0011100000100011    0011100000100100    0011100000100101    0011100000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14370 - 14374

  --0011100000100111    0011100000101000    0011100000101001    0011100000101010    0011100000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14375 - 14379

  --0011100000101100    0011100000101101    0011100000101110    0011100000101111    0011100000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14380 - 14384

  --0011100000110001    0011100000110010    0011100000110011    0011100000110100    0011100000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14385 - 14389

  --0011100000110110    0011100000110111    0011100000111000    0011100000111001    0011100000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14390 - 14394

  --0011100000111011    0011100000111100    0011100000111101    0011100000111110    0011100000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14395 - 14399

  --0011100001000000    0011100001000001    0011100001000010    0011100001000011    0011100001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14400 - 14404

  --0011100001000101    0011100001000110    0011100001000111    0011100001001000    0011100001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14405 - 14409

  --0011100001001010    0011100001001011    0011100001001100    0011100001001101    0011100001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14410 - 14414

  --0011100001001111    0011100001010000    0011100001010001    0011100001010010    0011100001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14415 - 14419

  --0011100001010100    0011100001010101    0011100001010110    0011100001010111    0011100001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14420 - 14424

  --0011100001011001    0011100001011010    0011100001011011    0011100001011100    0011100001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14425 - 14429

  --0011100001011110    0011100001011111    0011100001100000    0011100001100001    0011100001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14430 - 14434

  --0011100001100011    0011100001100100    0011100001100101    0011100001100110    0011100001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14435 - 14439

  --0011100001101000    0011100001101001    0011100001101010    0011100001101011    0011100001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14440 - 14444

  --0011100001101101    0011100001101110    0011100001101111    0011100001110000    0011100001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14445 - 14449

  --0011100001110010    0011100001110011    0011100001110100    0011100001110101    0011100001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14450 - 14454

  --0011100001110111    0011100001111000    0011100001111001    0011100001111010    0011100001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14455 - 14459

  --0011100001111100    0011100001111101    0011100001111110    0011100001111111    0011100010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14460 - 14464

  --0011100010000001    0011100010000010    0011100010000011    0011100010000100    0011100010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14465 - 14469

  --0011100010000110    0011100010000111    0011100010001000    0011100010001001    0011100010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14470 - 14474

  --0011100010001011    0011100010001100    0011100010001101    0011100010001110    0011100010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14475 - 14479

  --0011100010010000    0011100010010001    0011100010010010    0011100010010011    0011100010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14480 - 14484

  --0011100010010101    0011100010010110    0011100010010111    0011100010011000    0011100010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14485 - 14489

  --0011100010011010    0011100010011011    0011100010011100    0011100010011101    0011100010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14490 - 14494

  --0011100010011111    0011100010100000    0011100010100001    0011100010100010    0011100010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14495 - 14499

  --0011100010100100    0011100010100101    0011100010100110    0011100010100111    0011100010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14500 - 14504

  --0011100010101001    0011100010101010    0011100010101011    0011100010101100    0011100010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14505 - 14509

  --0011100010101110    0011100010101111    0011100010110000    0011100010110001    0011100010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14510 - 14514

  --0011100010110011    0011100010110100    0011100010110101    0011100010110110    0011100010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14515 - 14519

  --0011100010111000    0011100010111001    0011100010111010    0011100010111011    0011100010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14520 - 14524

  --0011100010111101    0011100010111110    0011100010111111    0011100011000000    0011100011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14525 - 14529

  --0011100011000010    0011100011000011    0011100011000100    0011100011000101    0011100011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14530 - 14534

  --0011100011000111    0011100011001000    0011100011001001    0011100011001010    0011100011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14535 - 14539

  --0011100011001100    0011100011001101    0011100011001110    0011100011001111    0011100011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14540 - 14544

  --0011100011010001    0011100011010010    0011100011010011    0011100011010100    0011100011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14545 - 14549

  --0011100011010110    0011100011010111    0011100011011000    0011100011011001    0011100011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14550 - 14554

  --0011100011011011    0011100011011100    0011100011011101    0011100011011110    0011100011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14555 - 14559

  --0011100011100000    0011100011100001    0011100011100010    0011100011100011    0011100011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14560 - 14564

  --0011100011100101    0011100011100110    0011100011100111    0011100011101000    0011100011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14565 - 14569

  --0011100011101010    0011100011101011    0011100011101100    0011100011101101    0011100011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14570 - 14574

  --0011100011101111    0011100011110000    0011100011110001    0011100011110010    0011100011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14575 - 14579

  --0011100011110100    0011100011110101    0011100011110110    0011100011110111    0011100011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14580 - 14584

  --0011100011111001    0011100011111010    0011100011111011    0011100011111100    0011100011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14585 - 14589

  --0011100011111110    0011100011111111    0011100100000000    0011100100000001    0011100100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14590 - 14594

  --0011100100000011    0011100100000100    0011100100000101    0011100100000110    0011100100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14595 - 14599

  --0011100100001000    0011100100001001    0011100100001010    0011100100001011    0011100100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14600 - 14604

  --0011100100001101    0011100100001110    0011100100001111    0011100100010000    0011100100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14605 - 14609

  --0011100100010010    0011100100010011    0011100100010100    0011100100010101    0011100100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14610 - 14614

  --0011100100010111    0011100100011000    0011100100011001    0011100100011010    0011100100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14615 - 14619

  --0011100100011100    0011100100011101    0011100100011110    0011100100011111    0011100100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14620 - 14624

  --0011100100100001    0011100100100010    0011100100100011    0011100100100100    0011100100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14625 - 14629

  --0011100100100110    0011100100100111    0011100100101000    0011100100101001    0011100100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14630 - 14634

  --0011100100101011    0011100100101100    0011100100101101    0011100100101110    0011100100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14635 - 14639

  --0011100100110000    0011100100110001    0011100100110010    0011100100110011    0011100100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14640 - 14644

  --0011100100110101    0011100100110110    0011100100110111    0011100100111000    0011100100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14645 - 14649

  --0011100100111010    0011100100111011    0011100100111100    0011100100111101    0011100100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14650 - 14654

  --0011100100111111    0011100101000000    0011100101000001    0011100101000010    0011100101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14655 - 14659

  --0011100101000100    0011100101000101    0011100101000110    0011100101000111    0011100101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14660 - 14664

  --0011100101001001    0011100101001010    0011100101001011    0011100101001100    0011100101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14665 - 14669

  --0011100101001110    0011100101001111    0011100101010000    0011100101010001    0011100101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14670 - 14674

  --0011100101010011    0011100101010100    0011100101010101    0011100101010110    0011100101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14675 - 14679

  --0011100101011000    0011100101011001    0011100101011010    0011100101011011    0011100101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14680 - 14684

  --0011100101011101    0011100101011110    0011100101011111    0011100101100000    0011100101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14685 - 14689

  --0011100101100010    0011100101100011    0011100101100100    0011100101100101    0011100101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14690 - 14694

  --0011100101100111    0011100101101000    0011100101101001    0011100101101010    0011100101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14695 - 14699

  --0011100101101100    0011100101101101    0011100101101110    0011100101101111    0011100101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14700 - 14704

  --0011100101110001    0011100101110010    0011100101110011    0011100101110100    0011100101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14705 - 14709

  --0011100101110110    0011100101110111    0011100101111000    0011100101111001    0011100101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14710 - 14714

  --0011100101111011    0011100101111100    0011100101111101    0011100101111110    0011100101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14715 - 14719

  --0011100110000000    0011100110000001    0011100110000010    0011100110000011    0011100110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14720 - 14724

  --0011100110000101    0011100110000110    0011100110000111    0011100110001000    0011100110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14725 - 14729

  --0011100110001010    0011100110001011    0011100110001100    0011100110001101    0011100110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14730 - 14734

  --0011100110001111    0011100110010000    0011100110010001    0011100110010010    0011100110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14735 - 14739

  --0011100110010100    0011100110010101    0011100110010110    0011100110010111    0011100110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14740 - 14744

  --0011100110011001    0011100110011010    0011100110011011    0011100110011100    0011100110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14745 - 14749

  --0011100110011110    0011100110011111    0011100110100000    0011100110100001    0011100110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14750 - 14754

  --0011100110100011    0011100110100100    0011100110100101    0011100110100110    0011100110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14755 - 14759

  --0011100110101000    0011100110101001    0011100110101010    0011100110101011    0011100110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14760 - 14764

  --0011100110101101    0011100110101110    0011100110101111    0011100110110000    0011100110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14765 - 14769

  --0011100110110010    0011100110110011    0011100110110100    0011100110110101    0011100110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14770 - 14774

  --0011100110110111    0011100110111000    0011100110111001    0011100110111010    0011100110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14775 - 14779

  --0011100110111100    0011100110111101    0011100110111110    0011100110111111    0011100111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14780 - 14784

  --0011100111000001    0011100111000010    0011100111000011    0011100111000100    0011100111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14785 - 14789

  --0011100111000110    0011100111000111    0011100111001000    0011100111001001    0011100111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14790 - 14794

  --0011100111001011    0011100111001100    0011100111001101    0011100111001110    0011100111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14795 - 14799

  --0011100111010000    0011100111010001    0011100111010010    0011100111010011    0011100111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14800 - 14804

  --0011100111010101    0011100111010110    0011100111010111    0011100111011000    0011100111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14805 - 14809

  --0011100111011010    0011100111011011    0011100111011100    0011100111011101    0011100111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14810 - 14814

  --0011100111011111    0011100111100000    0011100111100001    0011100111100010    0011100111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14815 - 14819

  --0011100111100100    0011100111100101    0011100111100110    0011100111100111    0011100111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14820 - 14824

  --0011100111101001    0011100111101010    0011100111101011    0011100111101100    0011100111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14825 - 14829

  --0011100111101110    0011100111101111    0011100111110000    0011100111110001    0011100111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14830 - 14834

  --0011100111110011    0011100111110100    0011100111110101    0011100111110110    0011100111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14835 - 14839

  --0011100111111000    0011100111111001    0011100111111010    0011100111111011    0011100111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14840 - 14844

  --0011100111111101    0011100111111110    0011100111111111    0011101000000000    0011101000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14845 - 14849

  --0011101000000010    0011101000000011    0011101000000100    0011101000000101    0011101000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14850 - 14854

  --0011101000000111    0011101000001000    0011101000001001    0011101000001010    0011101000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14855 - 14859

  --0011101000001100    0011101000001101    0011101000001110    0011101000001111    0011101000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14860 - 14864

  --0011101000010001    0011101000010010    0011101000010011    0011101000010100    0011101000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14865 - 14869

  --0011101000010110    0011101000010111    0011101000011000    0011101000011001    0011101000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14870 - 14874

  --0011101000011011    0011101000011100    0011101000011101    0011101000011110    0011101000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14875 - 14879

  --0011101000100000    0011101000100001    0011101000100010    0011101000100011    0011101000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14880 - 14884

  --0011101000100101    0011101000100110    0011101000100111    0011101000101000    0011101000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14885 - 14889

  --0011101000101010    0011101000101011    0011101000101100    0011101000101101    0011101000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14890 - 14894

  --0011101000101111    0011101000110000    0011101000110001    0011101000110010    0011101000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14895 - 14899

  --0011101000110100    0011101000110101    0011101000110110    0011101000110111    0011101000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14900 - 14904

  --0011101000111001    0011101000111010    0011101000111011    0011101000111100    0011101000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14905 - 14909

  --0011101000111110    0011101000111111    0011101001000000    0011101001000001    0011101001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14910 - 14914

  --0011101001000011    0011101001000100    0011101001000101    0011101001000110    0011101001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14915 - 14919

  --0011101001001000    0011101001001001    0011101001001010    0011101001001011    0011101001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14920 - 14924

  --0011101001001101    0011101001001110    0011101001001111    0011101001010000    0011101001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14925 - 14929

  --0011101001010010    0011101001010011    0011101001010100    0011101001010101    0011101001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14930 - 14934

  --0011101001010111    0011101001011000    0011101001011001    0011101001011010    0011101001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14935 - 14939

  --0011101001011100    0011101001011101    0011101001011110    0011101001011111    0011101001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14940 - 14944

  --0011101001100001    0011101001100010    0011101001100011    0011101001100100    0011101001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14945 - 14949

  --0011101001100110    0011101001100111    0011101001101000    0011101001101001    0011101001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14950 - 14954

  --0011101001101011    0011101001101100    0011101001101101    0011101001101110    0011101001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14955 - 14959

  --0011101001110000    0011101001110001    0011101001110010    0011101001110011    0011101001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14960 - 14964

  --0011101001110101    0011101001110110    0011101001110111    0011101001111000    0011101001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14965 - 14969

  --0011101001111010    0011101001111011    0011101001111100    0011101001111101    0011101001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14970 - 14974

  --0011101001111111    0011101010000000    0011101010000001    0011101010000010    0011101010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14975 - 14979

  --0011101010000100    0011101010000101    0011101010000110    0011101010000111    0011101010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14980 - 14984

  --0011101010001001    0011101010001010    0011101010001011    0011101010001100    0011101010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14985 - 14989

  --0011101010001110    0011101010001111    0011101010010000    0011101010010001    0011101010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14990 - 14994

  --0011101010010011    0011101010010100    0011101010010101    0011101010010110    0011101010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 14995 - 14999

  --0011101010011000    0011101010011001    0011101010011010    0011101010011011    0011101010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15000 - 15004

  --0011101010011101    0011101010011110    0011101010011111    0011101010100000    0011101010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15005 - 15009

  --0011101010100010    0011101010100011    0011101010100100    0011101010100101    0011101010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15010 - 15014

  --0011101010100111    0011101010101000    0011101010101001    0011101010101010    0011101010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15015 - 15019

  --0011101010101100    0011101010101101    0011101010101110    0011101010101111    0011101010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15020 - 15024

  --0011101010110001    0011101010110010    0011101010110011    0011101010110100    0011101010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15025 - 15029

  --0011101010110110    0011101010110111    0011101010111000    0011101010111001    0011101010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15030 - 15034

  --0011101010111011    0011101010111100    0011101010111101    0011101010111110    0011101010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15035 - 15039

  --0011101011000000    0011101011000001    0011101011000010    0011101011000011    0011101011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15040 - 15044

  --0011101011000101    0011101011000110    0011101011000111    0011101011001000    0011101011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15045 - 15049

  --0011101011001010    0011101011001011    0011101011001100    0011101011001101    0011101011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15050 - 15054

  --0011101011001111    0011101011010000    0011101011010001    0011101011010010    0011101011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15055 - 15059

  --0011101011010100    0011101011010101    0011101011010110    0011101011010111    0011101011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15060 - 15064

  --0011101011011001    0011101011011010    0011101011011011    0011101011011100    0011101011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15065 - 15069

  --0011101011011110    0011101011011111    0011101011100000    0011101011100001    0011101011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15070 - 15074

  --0011101011100011    0011101011100100    0011101011100101    0011101011100110    0011101011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15075 - 15079

  --0011101011101000    0011101011101001    0011101011101010    0011101011101011    0011101011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15080 - 15084

  --0011101011101101    0011101011101110    0011101011101111    0011101011110000    0011101011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15085 - 15089

  --0011101011110010    0011101011110011    0011101011110100    0011101011110101    0011101011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15090 - 15094

  --0011101011110111    0011101011111000    0011101011111001    0011101011111010    0011101011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15095 - 15099

  --0011101011111100    0011101011111101    0011101011111110    0011101011111111    0011101100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15100 - 15104

  --0011101100000001    0011101100000010    0011101100000011    0011101100000100    0011101100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15105 - 15109

  --0011101100000110    0011101100000111    0011101100001000    0011101100001001    0011101100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15110 - 15114

  --0011101100001011    0011101100001100    0011101100001101    0011101100001110    0011101100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15115 - 15119

  --0011101100010000    0011101100010001    0011101100010010    0011101100010011    0011101100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15120 - 15124

  --0011101100010101    0011101100010110    0011101100010111    0011101100011000    0011101100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15125 - 15129

  --0011101100011010    0011101100011011    0011101100011100    0011101100011101    0011101100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15130 - 15134

  --0011101100011111    0011101100100000    0011101100100001    0011101100100010    0011101100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15135 - 15139

  --0011101100100100    0011101100100101    0011101100100110    0011101100100111    0011101100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15140 - 15144

  --0011101100101001    0011101100101010    0011101100101011    0011101100101100    0011101100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15145 - 15149

  --0011101100101110    0011101100101111    0011101100110000    0011101100110001    0011101100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15150 - 15154

  --0011101100110011    0011101100110100    0011101100110101    0011101100110110    0011101100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15155 - 15159

  --0011101100111000    0011101100111001    0011101100111010    0011101100111011    0011101100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15160 - 15164

  --0011101100111101    0011101100111110    0011101100111111    0011101101000000    0011101101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15165 - 15169

  --0011101101000010    0011101101000011    0011101101000100    0011101101000101    0011101101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15170 - 15174

  --0011101101000111    0011101101001000    0011101101001001    0011101101001010    0011101101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15175 - 15179

  --0011101101001100    0011101101001101    0011101101001110    0011101101001111    0011101101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15180 - 15184

  --0011101101010001    0011101101010010    0011101101010011    0011101101010100    0011101101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15185 - 15189

  --0011101101010110    0011101101010111    0011101101011000    0011101101011001    0011101101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15190 - 15194

  --0011101101011011    0011101101011100    0011101101011101    0011101101011110    0011101101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15195 - 15199

  --0011101101100000    0011101101100001    0011101101100010    0011101101100011    0011101101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15200 - 15204

  --0011101101100101    0011101101100110    0011101101100111    0011101101101000    0011101101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15205 - 15209

  --0011101101101010    0011101101101011    0011101101101100    0011101101101101    0011101101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15210 - 15214

  --0011101101101111    0011101101110000    0011101101110001    0011101101110010    0011101101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15215 - 15219

  --0011101101110100    0011101101110101    0011101101110110    0011101101110111    0011101101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15220 - 15224

  --0011101101111001    0011101101111010    0011101101111011    0011101101111100    0011101101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15225 - 15229

  --0011101101111110    0011101101111111    0011101110000000    0011101110000001    0011101110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15230 - 15234

  --0011101110000011    0011101110000100    0011101110000101    0011101110000110    0011101110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15235 - 15239

  --0011101110001000    0011101110001001    0011101110001010    0011101110001011    0011101110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15240 - 15244

  --0011101110001101    0011101110001110    0011101110001111    0011101110010000    0011101110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15245 - 15249

  --0011101110010010    0011101110010011    0011101110010100    0011101110010101    0011101110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15250 - 15254

  --0011101110010111    0011101110011000    0011101110011001    0011101110011010    0011101110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15255 - 15259

  --0011101110011100    0011101110011101    0011101110011110    0011101110011111    0011101110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15260 - 15264

  --0011101110100001    0011101110100010    0011101110100011    0011101110100100    0011101110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15265 - 15269

  --0011101110100110    0011101110100111    0011101110101000    0011101110101001    0011101110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15270 - 15274

  --0011101110101011    0011101110101100    0011101110101101    0011101110101110    0011101110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15275 - 15279

  --0011101110110000    0011101110110001    0011101110110010    0011101110110011    0011101110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15280 - 15284

  --0011101110110101    0011101110110110    0011101110110111    0011101110111000    0011101110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15285 - 15289

  --0011101110111010    0011101110111011    0011101110111100    0011101110111101    0011101110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15290 - 15294

  --0011101110111111    0011101111000000    0011101111000001    0011101111000010    0011101111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15295 - 15299

  --0011101111000100    0011101111000101    0011101111000110    0011101111000111    0011101111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15300 - 15304

  --0011101111001001    0011101111001010    0011101111001011    0011101111001100    0011101111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15305 - 15309

  --0011101111001110    0011101111001111    0011101111010000    0011101111010001    0011101111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15310 - 15314

  --0011101111010011    0011101111010100    0011101111010101    0011101111010110    0011101111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15315 - 15319

  --0011101111011000    0011101111011001    0011101111011010    0011101111011011    0011101111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15320 - 15324

  --0011101111011101    0011101111011110    0011101111011111    0011101111100000    0011101111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15325 - 15329

  --0011101111100010    0011101111100011    0011101111100100    0011101111100101    0011101111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15330 - 15334

  --0011101111100111    0011101111101000    0011101111101001    0011101111101010    0011101111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15335 - 15339

  --0011101111101100    0011101111101101    0011101111101110    0011101111101111    0011101111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15340 - 15344

  --0011101111110001    0011101111110010    0011101111110011    0011101111110100    0011101111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15345 - 15349

  --0011101111110110    0011101111110111    0011101111111000    0011101111111001    0011101111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15350 - 15354

  --0011101111111011    0011101111111100    0011101111111101    0011101111111110    0011101111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15355 - 15359

  --0011110000000000    0011110000000001    0011110000000010    0011110000000011    0011110000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15360 - 15364

  --0011110000000101    0011110000000110    0011110000000111    0011110000001000    0011110000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15365 - 15369

  --0011110000001010    0011110000001011    0011110000001100    0011110000001101    0011110000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15370 - 15374

  --0011110000001111    0011110000010000    0011110000010001    0011110000010010    0011110000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15375 - 15379

  --0011110000010100    0011110000010101    0011110000010110    0011110000010111    0011110000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15380 - 15384

  --0011110000011001    0011110000011010    0011110000011011    0011110000011100    0011110000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15385 - 15389

  --0011110000011110    0011110000011111    0011110000100000    0011110000100001    0011110000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15390 - 15394

  --0011110000100011    0011110000100100    0011110000100101    0011110000100110    0011110000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15395 - 15399

  --0011110000101000    0011110000101001    0011110000101010    0011110000101011    0011110000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15400 - 15404

  --0011110000101101    0011110000101110    0011110000101111    0011110000110000    0011110000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15405 - 15409

  --0011110000110010    0011110000110011    0011110000110100    0011110000110101    0011110000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15410 - 15414

  --0011110000110111    0011110000111000    0011110000111001    0011110000111010    0011110000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15415 - 15419

  --0011110000111100    0011110000111101    0011110000111110    0011110000111111    0011110001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15420 - 15424

  --0011110001000001    0011110001000010    0011110001000011    0011110001000100    0011110001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15425 - 15429

  --0011110001000110    0011110001000111    0011110001001000    0011110001001001    0011110001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15430 - 15434

  --0011110001001011    0011110001001100    0011110001001101    0011110001001110    0011110001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15435 - 15439

  --0011110001010000    0011110001010001    0011110001010010    0011110001010011    0011110001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15440 - 15444

  --0011110001010101    0011110001010110    0011110001010111    0011110001011000    0011110001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15445 - 15449

  --0011110001011010    0011110001011011    0011110001011100    0011110001011101    0011110001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15450 - 15454

  --0011110001011111    0011110001100000    0011110001100001    0011110001100010    0011110001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15455 - 15459

  --0011110001100100    0011110001100101    0011110001100110    0011110001100111    0011110001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15460 - 15464

  --0011110001101001    0011110001101010    0011110001101011    0011110001101100    0011110001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15465 - 15469

  --0011110001101110    0011110001101111    0011110001110000    0011110001110001    0011110001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15470 - 15474

  --0011110001110011    0011110001110100    0011110001110101    0011110001110110    0011110001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15475 - 15479

  --0011110001111000    0011110001111001    0011110001111010    0011110001111011    0011110001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15480 - 15484

  --0011110001111101    0011110001111110    0011110001111111    0011110010000000    0011110010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15485 - 15489

  --0011110010000010    0011110010000011    0011110010000100    0011110010000101    0011110010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15490 - 15494

  --0011110010000111    0011110010001000    0011110010001001    0011110010001010    0011110010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15495 - 15499

  --0011110010001100    0011110010001101    0011110010001110    0011110010001111    0011110010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15500 - 15504

  --0011110010010001    0011110010010010    0011110010010011    0011110010010100    0011110010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15505 - 15509

  --0011110010010110    0011110010010111    0011110010011000    0011110010011001    0011110010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15510 - 15514

  --0011110010011011    0011110010011100    0011110010011101    0011110010011110    0011110010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15515 - 15519

  --0011110010100000    0011110010100001    0011110010100010    0011110010100011    0011110010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15520 - 15524

  --0011110010100101    0011110010100110    0011110010100111    0011110010101000    0011110010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15525 - 15529

  --0011110010101010    0011110010101011    0011110010101100    0011110010101101    0011110010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15530 - 15534

  --0011110010101111    0011110010110000    0011110010110001    0011110010110010    0011110010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15535 - 15539

  --0011110010110100    0011110010110101    0011110010110110    0011110010110111    0011110010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15540 - 15544

  --0011110010111001    0011110010111010    0011110010111011    0011110010111100    0011110010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15545 - 15549

  --0011110010111110    0011110010111111    0011110011000000    0011110011000001    0011110011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15550 - 15554

  --0011110011000011    0011110011000100    0011110011000101    0011110011000110    0011110011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15555 - 15559

  --0011110011001000    0011110011001001    0011110011001010    0011110011001011    0011110011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15560 - 15564

  --0011110011001101    0011110011001110    0011110011001111    0011110011010000    0011110011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15565 - 15569

  --0011110011010010    0011110011010011    0011110011010100    0011110011010101    0011110011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15570 - 15574

  --0011110011010111    0011110011011000    0011110011011001    0011110011011010    0011110011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15575 - 15579

  --0011110011011100    0011110011011101    0011110011011110    0011110011011111    0011110011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15580 - 15584

  --0011110011100001    0011110011100010    0011110011100011    0011110011100100    0011110011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15585 - 15589

  --0011110011100110    0011110011100111    0011110011101000    0011110011101001    0011110011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15590 - 15594

  --0011110011101011    0011110011101100    0011110011101101    0011110011101110    0011110011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15595 - 15599

  --0011110011110000    0011110011110001    0011110011110010    0011110011110011    0011110011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15600 - 15604

  --0011110011110101    0011110011110110    0011110011110111    0011110011111000    0011110011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15605 - 15609

  --0011110011111010    0011110011111011    0011110011111100    0011110011111101    0011110011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15610 - 15614

  --0011110011111111    0011110100000000    0011110100000001    0011110100000010    0011110100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15615 - 15619

  --0011110100000100    0011110100000101    0011110100000110    0011110100000111    0011110100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15620 - 15624

  --0011110100001001    0011110100001010    0011110100001011    0011110100001100    0011110100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15625 - 15629

  --0011110100001110    0011110100001111    0011110100010000    0011110100010001    0011110100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15630 - 15634

  --0011110100010011    0011110100010100    0011110100010101    0011110100010110    0011110100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15635 - 15639

  --0011110100011000    0011110100011001    0011110100011010    0011110100011011    0011110100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15640 - 15644

  --0011110100011101    0011110100011110    0011110100011111    0011110100100000    0011110100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15645 - 15649

  --0011110100100010    0011110100100011    0011110100100100    0011110100100101    0011110100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15650 - 15654

  --0011110100100111    0011110100101000    0011110100101001    0011110100101010    0011110100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15655 - 15659

  --0011110100101100    0011110100101101    0011110100101110    0011110100101111    0011110100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15660 - 15664

  --0011110100110001    0011110100110010    0011110100110011    0011110100110100    0011110100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15665 - 15669

  --0011110100110110    0011110100110111    0011110100111000    0011110100111001    0011110100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15670 - 15674

  --0011110100111011    0011110100111100    0011110100111101    0011110100111110    0011110100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15675 - 15679

  --0011110101000000    0011110101000001    0011110101000010    0011110101000011    0011110101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15680 - 15684

  --0011110101000101    0011110101000110    0011110101000111    0011110101001000    0011110101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15685 - 15689

  --0011110101001010    0011110101001011    0011110101001100    0011110101001101    0011110101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15690 - 15694

  --0011110101001111    0011110101010000    0011110101010001    0011110101010010    0011110101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15695 - 15699

  --0011110101010100    0011110101010101    0011110101010110    0011110101010111    0011110101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15700 - 15704

  --0011110101011001    0011110101011010    0011110101011011    0011110101011100    0011110101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15705 - 15709

  --0011110101011110    0011110101011111    0011110101100000    0011110101100001    0011110101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15710 - 15714

  --0011110101100011    0011110101100100    0011110101100101    0011110101100110    0011110101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15715 - 15719

  --0011110101101000    0011110101101001    0011110101101010    0011110101101011    0011110101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15720 - 15724

  --0011110101101101    0011110101101110    0011110101101111    0011110101110000    0011110101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15725 - 15729

  --0011110101110010    0011110101110011    0011110101110100    0011110101110101    0011110101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15730 - 15734

  --0011110101110111    0011110101111000    0011110101111001    0011110101111010    0011110101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15735 - 15739

  --0011110101111100    0011110101111101    0011110101111110    0011110101111111    0011110110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15740 - 15744

  --0011110110000001    0011110110000010    0011110110000011    0011110110000100    0011110110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15745 - 15749

  --0011110110000110    0011110110000111    0011110110001000    0011110110001001    0011110110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15750 - 15754

  --0011110110001011    0011110110001100    0011110110001101    0011110110001110    0011110110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15755 - 15759

  --0011110110010000    0011110110010001    0011110110010010    0011110110010011    0011110110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15760 - 15764

  --0011110110010101    0011110110010110    0011110110010111    0011110110011000    0011110110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15765 - 15769

  --0011110110011010    0011110110011011    0011110110011100    0011110110011101    0011110110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15770 - 15774

  --0011110110011111    0011110110100000    0011110110100001    0011110110100010    0011110110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15775 - 15779

  --0011110110100100    0011110110100101    0011110110100110    0011110110100111    0011110110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15780 - 15784

  --0011110110101001    0011110110101010    0011110110101011    0011110110101100    0011110110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15785 - 15789

  --0011110110101110    0011110110101111    0011110110110000    0011110110110001    0011110110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15790 - 15794

  --0011110110110011    0011110110110100    0011110110110101    0011110110110110    0011110110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15795 - 15799

  --0011110110111000    0011110110111001    0011110110111010    0011110110111011    0011110110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15800 - 15804

  --0011110110111101    0011110110111110    0011110110111111    0011110111000000    0011110111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15805 - 15809

  --0011110111000010    0011110111000011    0011110111000100    0011110111000101    0011110111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15810 - 15814

  --0011110111000111    0011110111001000    0011110111001001    0011110111001010    0011110111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15815 - 15819

  --0011110111001100    0011110111001101    0011110111001110    0011110111001111    0011110111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15820 - 15824

  --0011110111010001    0011110111010010    0011110111010011    0011110111010100    0011110111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15825 - 15829

  --0011110111010110    0011110111010111    0011110111011000    0011110111011001    0011110111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15830 - 15834

  --0011110111011011    0011110111011100    0011110111011101    0011110111011110    0011110111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15835 - 15839

  --0011110111100000    0011110111100001    0011110111100010    0011110111100011    0011110111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15840 - 15844

  --0011110111100101    0011110111100110    0011110111100111    0011110111101000    0011110111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15845 - 15849

  --0011110111101010    0011110111101011    0011110111101100    0011110111101101    0011110111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15850 - 15854

  --0011110111101111    0011110111110000    0011110111110001    0011110111110010    0011110111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15855 - 15859

  --0011110111110100    0011110111110101    0011110111110110    0011110111110111    0011110111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15860 - 15864

  --0011110111111001    0011110111111010    0011110111111011    0011110111111100    0011110111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15865 - 15869

  --0011110111111110    0011110111111111    0011111000000000    0011111000000001    0011111000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15870 - 15874

  --0011111000000011    0011111000000100    0011111000000101    0011111000000110    0011111000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15875 - 15879

  --0011111000001000    0011111000001001    0011111000001010    0011111000001011    0011111000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15880 - 15884

  --0011111000001101    0011111000001110    0011111000001111    0011111000010000    0011111000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15885 - 15889

  --0011111000010010    0011111000010011    0011111000010100    0011111000010101    0011111000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15890 - 15894

  --0011111000010111    0011111000011000    0011111000011001    0011111000011010    0011111000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15895 - 15899

  --0011111000011100    0011111000011101    0011111000011110    0011111000011111    0011111000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15900 - 15904

  --0011111000100001    0011111000100010    0011111000100011    0011111000100100    0011111000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15905 - 15909

  --0011111000100110    0011111000100111    0011111000101000    0011111000101001    0011111000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15910 - 15914

  --0011111000101011    0011111000101100    0011111000101101    0011111000101110    0011111000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15915 - 15919

  --0011111000110000    0011111000110001    0011111000110010    0011111000110011    0011111000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15920 - 15924

  --0011111000110101    0011111000110110    0011111000110111    0011111000111000    0011111000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15925 - 15929

  --0011111000111010    0011111000111011    0011111000111100    0011111000111101    0011111000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15930 - 15934

  --0011111000111111    0011111001000000    0011111001000001    0011111001000010    0011111001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15935 - 15939

  --0011111001000100    0011111001000101    0011111001000110    0011111001000111    0011111001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15940 - 15944

  --0011111001001001    0011111001001010    0011111001001011    0011111001001100    0011111001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15945 - 15949

  --0011111001001110    0011111001001111    0011111001010000    0011111001010001    0011111001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15950 - 15954

  --0011111001010011    0011111001010100    0011111001010101    0011111001010110    0011111001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15955 - 15959

  --0011111001011000    0011111001011001    0011111001011010    0011111001011011    0011111001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15960 - 15964

  --0011111001011101    0011111001011110    0011111001011111    0011111001100000    0011111001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15965 - 15969

  --0011111001100010    0011111001100011    0011111001100100    0011111001100101    0011111001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15970 - 15974

  --0011111001100111    0011111001101000    0011111001101001    0011111001101010    0011111001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15975 - 15979

  --0011111001101100    0011111001101101    0011111001101110    0011111001101111    0011111001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15980 - 15984

  --0011111001110001    0011111001110010    0011111001110011    0011111001110100    0011111001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15985 - 15989

  --0011111001110110    0011111001110111    0011111001111000    0011111001111001    0011111001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15990 - 15994

  --0011111001111011    0011111001111100    0011111001111101    0011111001111110    0011111001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 15995 - 15999

  --0011111010000000    0011111010000001    0011111010000010    0011111010000011    0011111010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16000 - 16004

  --0011111010000101    0011111010000110    0011111010000111    0011111010001000    0011111010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16005 - 16009

  --0011111010001010    0011111010001011    0011111010001100    0011111010001101    0011111010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16010 - 16014

  --0011111010001111    0011111010010000    0011111010010001    0011111010010010    0011111010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16015 - 16019

  --0011111010010100    0011111010010101    0011111010010110    0011111010010111    0011111010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16020 - 16024

  --0011111010011001    0011111010011010    0011111010011011    0011111010011100    0011111010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16025 - 16029

  --0011111010011110    0011111010011111    0011111010100000    0011111010100001    0011111010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16030 - 16034

  --0011111010100011    0011111010100100    0011111010100101    0011111010100110    0011111010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16035 - 16039

  --0011111010101000    0011111010101001    0011111010101010    0011111010101011    0011111010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16040 - 16044

  --0011111010101101    0011111010101110    0011111010101111    0011111010110000    0011111010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16045 - 16049

  --0011111010110010    0011111010110011    0011111010110100    0011111010110101    0011111010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16050 - 16054

  --0011111010110111    0011111010111000    0011111010111001    0011111010111010    0011111010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16055 - 16059

  --0011111010111100    0011111010111101    0011111010111110    0011111010111111    0011111011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16060 - 16064

  --0011111011000001    0011111011000010    0011111011000011    0011111011000100    0011111011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16065 - 16069

  --0011111011000110    0011111011000111    0011111011001000    0011111011001001    0011111011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16070 - 16074

  --0011111011001011    0011111011001100    0011111011001101    0011111011001110    0011111011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16075 - 16079

  --0011111011010000    0011111011010001    0011111011010010    0011111011010011    0011111011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16080 - 16084

  --0011111011010101    0011111011010110    0011111011010111    0011111011011000    0011111011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16085 - 16089

  --0011111011011010    0011111011011011    0011111011011100    0011111011011101    0011111011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16090 - 16094

  --0011111011011111    0011111011100000    0011111011100001    0011111011100010    0011111011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16095 - 16099

  --0011111011100100    0011111011100101    0011111011100110    0011111011100111    0011111011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16100 - 16104

  --0011111011101001    0011111011101010    0011111011101011    0011111011101100    0011111011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16105 - 16109

  --0011111011101110    0011111011101111    0011111011110000    0011111011110001    0011111011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16110 - 16114

  --0011111011110011    0011111011110100    0011111011110101    0011111011110110    0011111011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16115 - 16119

  --0011111011111000    0011111011111001    0011111011111010    0011111011111011    0011111011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16120 - 16124

  --0011111011111101    0011111011111110    0011111011111111    0011111100000000    0011111100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16125 - 16129

  --0011111100000010    0011111100000011    0011111100000100    0011111100000101    0011111100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16130 - 16134

  --0011111100000111    0011111100001000    0011111100001001    0011111100001010    0011111100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16135 - 16139

  --0011111100001100    0011111100001101    0011111100001110    0011111100001111    0011111100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16140 - 16144

  --0011111100010001    0011111100010010    0011111100010011    0011111100010100    0011111100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16145 - 16149

  --0011111100010110    0011111100010111    0011111100011000    0011111100011001    0011111100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16150 - 16154

  --0011111100011011    0011111100011100    0011111100011101    0011111100011110    0011111100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16155 - 16159

  --0011111100100000    0011111100100001    0011111100100010    0011111100100011    0011111100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16160 - 16164

  --0011111100100101    0011111100100110    0011111100100111    0011111100101000    0011111100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16165 - 16169

  --0011111100101010    0011111100101011    0011111100101100    0011111100101101    0011111100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16170 - 16174

  --0011111100101111    0011111100110000    0011111100110001    0011111100110010    0011111100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16175 - 16179

  --0011111100110100    0011111100110101    0011111100110110    0011111100110111    0011111100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16180 - 16184

  --0011111100111001    0011111100111010    0011111100111011    0011111100111100    0011111100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16185 - 16189

  --0011111100111110    0011111100111111    0011111101000000    0011111101000001    0011111101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16190 - 16194

  --0011111101000011    0011111101000100    0011111101000101    0011111101000110    0011111101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16195 - 16199

  --0011111101001000    0011111101001001    0011111101001010    0011111101001011    0011111101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16200 - 16204

  --0011111101001101    0011111101001110    0011111101001111    0011111101010000    0011111101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16205 - 16209

  --0011111101010010    0011111101010011    0011111101010100    0011111101010101    0011111101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16210 - 16214

  --0011111101010111    0011111101011000    0011111101011001    0011111101011010    0011111101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16215 - 16219

  --0011111101011100    0011111101011101    0011111101011110    0011111101011111    0011111101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16220 - 16224

  --0011111101100001    0011111101100010    0011111101100011    0011111101100100    0011111101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16225 - 16229

  --0011111101100110    0011111101100111    0011111101101000    0011111101101001    0011111101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16230 - 16234

  --0011111101101011    0011111101101100    0011111101101101    0011111101101110    0011111101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16235 - 16239

  --0011111101110000    0011111101110001    0011111101110010    0011111101110011    0011111101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16240 - 16244

  --0011111101110101    0011111101110110    0011111101110111    0011111101111000    0011111101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16245 - 16249

  --0011111101111010    0011111101111011    0011111101111100    0011111101111101    0011111101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16250 - 16254

  --0011111101111111    0011111110000000    0011111110000001    0011111110000010    0011111110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16255 - 16259

  --0011111110000100    0011111110000101    0011111110000110    0011111110000111    0011111110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16260 - 16264

  --0011111110001001    0011111110001010    0011111110001011    0011111110001100    0011111110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16265 - 16269

  --0011111110001110    0011111110001111    0011111110010000    0011111110010001    0011111110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16270 - 16274

  --0011111110010011    0011111110010100    0011111110010101    0011111110010110    0011111110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16275 - 16279

  --0011111110011000    0011111110011001    0011111110011010    0011111110011011    0011111110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16280 - 16284

  --0011111110011101    0011111110011110    0011111110011111    0011111110100000    0011111110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16285 - 16289

  --0011111110100010    0011111110100011    0011111110100100    0011111110100101    0011111110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16290 - 16294

  --0011111110100111    0011111110101000    0011111110101001    0011111110101010    0011111110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16295 - 16299

  --0011111110101100    0011111110101101    0011111110101110    0011111110101111    0011111110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16300 - 16304

  --0011111110110001    0011111110110010    0011111110110011    0011111110110100    0011111110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16305 - 16309

  --0011111110110110    0011111110110111    0011111110111000    0011111110111001    0011111110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16310 - 16314

  --0011111110111011    0011111110111100    0011111110111101    0011111110111110    0011111110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16315 - 16319

  --0011111111000000    0011111111000001    0011111111000010    0011111111000011    0011111111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16320 - 16324

  --0011111111000101    0011111111000110    0011111111000111    0011111111001000    0011111111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16325 - 16329

  --0011111111001010    0011111111001011    0011111111001100    0011111111001101    0011111111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16330 - 16334

  --0011111111001111    0011111111010000    0011111111010001    0011111111010010    0011111111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16335 - 16339

  --0011111111010100    0011111111010101    0011111111010110    0011111111010111    0011111111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16340 - 16344

  --0011111111011001    0011111111011010    0011111111011011    0011111111011100    0011111111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16345 - 16349

  --0011111111011110    0011111111011111    0011111111100000    0011111111100001    0011111111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16350 - 16354

  --0011111111100011    0011111111100100    0011111111100101    0011111111100110    0011111111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16355 - 16359

  --0011111111101000    0011111111101001    0011111111101010    0011111111101011    0011111111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16360 - 16364

  --0011111111101101    0011111111101110    0011111111101111    0011111111110000    0011111111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16365 - 16369

  --0011111111110010    0011111111110011    0011111111110100    0011111111110101    0011111111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16370 - 16374

  --0011111111110111    0011111111111000    0011111111111001    0011111111111010    0011111111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16375 - 16379

  --0011111111111100    0011111111111101    0011111111111110    0011111111111111    0100000000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16380 - 16384

  --0100000000000001    0100000000000010    0100000000000011    0100000000000100    0100000000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16385 - 16389

  --0100000000000110    0100000000000111    0100000000001000    0100000000001001    0100000000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16390 - 16394

  --0100000000001011    0100000000001100    0100000000001101    0100000000001110    0100000000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16395 - 16399

  --0100000000010000    0100000000010001    0100000000010010    0100000000010011    0100000000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16400 - 16404

  --0100000000010101    0100000000010110    0100000000010111    0100000000011000    0100000000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16405 - 16409

  --0100000000011010    0100000000011011    0100000000011100    0100000000011101    0100000000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16410 - 16414

  --0100000000011111    0100000000100000    0100000000100001    0100000000100010    0100000000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16415 - 16419

  --0100000000100100    0100000000100101    0100000000100110    0100000000100111    0100000000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16420 - 16424

  --0100000000101001    0100000000101010    0100000000101011    0100000000101100    0100000000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16425 - 16429

  --0100000000101110    0100000000101111    0100000000110000    0100000000110001    0100000000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16430 - 16434

  --0100000000110011    0100000000110100    0100000000110101    0100000000110110    0100000000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16435 - 16439

  --0100000000111000    0100000000111001    0100000000111010    0100000000111011    0100000000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16440 - 16444

  --0100000000111101    0100000000111110    0100000000111111    0100000001000000    0100000001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16445 - 16449

  --0100000001000010    0100000001000011    0100000001000100    0100000001000101    0100000001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16450 - 16454

  --0100000001000111    0100000001001000    0100000001001001    0100000001001010    0100000001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16455 - 16459

  --0100000001001100    0100000001001101    0100000001001110    0100000001001111    0100000001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16460 - 16464

  --0100000001010001    0100000001010010    0100000001010011    0100000001010100    0100000001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16465 - 16469

  --0100000001010110    0100000001010111    0100000001011000    0100000001011001    0100000001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16470 - 16474

  --0100000001011011    0100000001011100    0100000001011101    0100000001011110    0100000001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16475 - 16479

  --0100000001100000    0100000001100001    0100000001100010    0100000001100011    0100000001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16480 - 16484

  --0100000001100101    0100000001100110    0100000001100111    0100000001101000    0100000001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16485 - 16489

  --0100000001101010    0100000001101011    0100000001101100    0100000001101101    0100000001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16490 - 16494

  --0100000001101111    0100000001110000    0100000001110001    0100000001110010    0100000001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16495 - 16499

  --0100000001110100    0100000001110101    0100000001110110    0100000001110111    0100000001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16500 - 16504

  --0100000001111001    0100000001111010    0100000001111011    0100000001111100    0100000001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16505 - 16509

  --0100000001111110    0100000001111111    0100000010000000    0100000010000001    0100000010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16510 - 16514

  --0100000010000011    0100000010000100    0100000010000101    0100000010000110    0100000010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16515 - 16519

  --0100000010001000    0100000010001001    0100000010001010    0100000010001011    0100000010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16520 - 16524

  --0100000010001101    0100000010001110    0100000010001111    0100000010010000    0100000010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16525 - 16529

  --0100000010010010    0100000010010011    0100000010010100    0100000010010101    0100000010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16530 - 16534

  --0100000010010111    0100000010011000    0100000010011001    0100000010011010    0100000010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16535 - 16539

  --0100000010011100    0100000010011101    0100000010011110    0100000010011111    0100000010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16540 - 16544

  --0100000010100001    0100000010100010    0100000010100011    0100000010100100    0100000010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16545 - 16549

  --0100000010100110    0100000010100111    0100000010101000    0100000010101001    0100000010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16550 - 16554

  --0100000010101011    0100000010101100    0100000010101101    0100000010101110    0100000010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16555 - 16559

  --0100000010110000    0100000010110001    0100000010110010    0100000010110011    0100000010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16560 - 16564

  --0100000010110101    0100000010110110    0100000010110111    0100000010111000    0100000010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16565 - 16569

  --0100000010111010    0100000010111011    0100000010111100    0100000010111101    0100000010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16570 - 16574

  --0100000010111111    0100000011000000    0100000011000001    0100000011000010    0100000011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16575 - 16579

  --0100000011000100    0100000011000101    0100000011000110    0100000011000111    0100000011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16580 - 16584

  --0100000011001001    0100000011001010    0100000011001011    0100000011001100    0100000011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16585 - 16589

  --0100000011001110    0100000011001111    0100000011010000    0100000011010001    0100000011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16590 - 16594

  --0100000011010011    0100000011010100    0100000011010101    0100000011010110    0100000011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16595 - 16599

  --0100000011011000    0100000011011001    0100000011011010    0100000011011011    0100000011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16600 - 16604

  --0100000011011101    0100000011011110    0100000011011111    0100000011100000    0100000011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16605 - 16609

  --0100000011100010    0100000011100011    0100000011100100    0100000011100101    0100000011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16610 - 16614

  --0100000011100111    0100000011101000    0100000011101001    0100000011101010    0100000011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16615 - 16619

  --0100000011101100    0100000011101101    0100000011101110    0100000011101111    0100000011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16620 - 16624

  --0100000011110001    0100000011110010    0100000011110011    0100000011110100    0100000011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16625 - 16629

  --0100000011110110    0100000011110111    0100000011111000    0100000011111001    0100000011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16630 - 16634

  --0100000011111011    0100000011111100    0100000011111101    0100000011111110    0100000011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16635 - 16639

  --0100000100000000    0100000100000001    0100000100000010    0100000100000011    0100000100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16640 - 16644

  --0100000100000101    0100000100000110    0100000100000111    0100000100001000    0100000100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16645 - 16649

  --0100000100001010    0100000100001011    0100000100001100    0100000100001101    0100000100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16650 - 16654

  --0100000100001111    0100000100010000    0100000100010001    0100000100010010    0100000100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16655 - 16659

  --0100000100010100    0100000100010101    0100000100010110    0100000100010111    0100000100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16660 - 16664

  --0100000100011001    0100000100011010    0100000100011011    0100000100011100    0100000100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16665 - 16669

  --0100000100011110    0100000100011111    0100000100100000    0100000100100001    0100000100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16670 - 16674

  --0100000100100011    0100000100100100    0100000100100101    0100000100100110    0100000100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16675 - 16679

  --0100000100101000    0100000100101001    0100000100101010    0100000100101011    0100000100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16680 - 16684

  --0100000100101101    0100000100101110    0100000100101111    0100000100110000    0100000100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16685 - 16689

  --0100000100110010    0100000100110011    0100000100110100    0100000100110101    0100000100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16690 - 16694

  --0100000100110111    0100000100111000    0100000100111001    0100000100111010    0100000100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16695 - 16699

  --0100000100111100    0100000100111101    0100000100111110    0100000100111111    0100000101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16700 - 16704

  --0100000101000001    0100000101000010    0100000101000011    0100000101000100    0100000101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16705 - 16709

  --0100000101000110    0100000101000111    0100000101001000    0100000101001001    0100000101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16710 - 16714

  --0100000101001011    0100000101001100    0100000101001101    0100000101001110    0100000101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16715 - 16719

  --0100000101010000    0100000101010001    0100000101010010    0100000101010011    0100000101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16720 - 16724

  --0100000101010101    0100000101010110    0100000101010111    0100000101011000    0100000101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16725 - 16729

  --0100000101011010    0100000101011011    0100000101011100    0100000101011101    0100000101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16730 - 16734

  --0100000101011111    0100000101100000    0100000101100001    0100000101100010    0100000101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16735 - 16739

  --0100000101100100    0100000101100101    0100000101100110    0100000101100111    0100000101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16740 - 16744

  --0100000101101001    0100000101101010    0100000101101011    0100000101101100    0100000101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16745 - 16749

  --0100000101101110    0100000101101111    0100000101110000    0100000101110001    0100000101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16750 - 16754

  --0100000101110011    0100000101110100    0100000101110101    0100000101110110    0100000101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16755 - 16759

  --0100000101111000    0100000101111001    0100000101111010    0100000101111011    0100000101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16760 - 16764

  --0100000101111101    0100000101111110    0100000101111111    0100000110000000    0100000110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16765 - 16769

  --0100000110000010    0100000110000011    0100000110000100    0100000110000101    0100000110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16770 - 16774

  --0100000110000111    0100000110001000    0100000110001001    0100000110001010    0100000110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16775 - 16779

  --0100000110001100    0100000110001101    0100000110001110    0100000110001111    0100000110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16780 - 16784

  --0100000110010001    0100000110010010    0100000110010011    0100000110010100    0100000110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16785 - 16789

  --0100000110010110    0100000110010111    0100000110011000    0100000110011001    0100000110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16790 - 16794

  --0100000110011011    0100000110011100    0100000110011101    0100000110011110    0100000110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16795 - 16799

  --0100000110100000    0100000110100001    0100000110100010    0100000110100011    0100000110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16800 - 16804

  --0100000110100101    0100000110100110    0100000110100111    0100000110101000    0100000110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16805 - 16809

  --0100000110101010    0100000110101011    0100000110101100    0100000110101101    0100000110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16810 - 16814

  --0100000110101111    0100000110110000    0100000110110001    0100000110110010    0100000110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16815 - 16819

  --0100000110110100    0100000110110101    0100000110110110    0100000110110111    0100000110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16820 - 16824

  --0100000110111001    0100000110111010    0100000110111011    0100000110111100    0100000110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16825 - 16829

  --0100000110111110    0100000110111111    0100000111000000    0100000111000001    0100000111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16830 - 16834

  --0100000111000011    0100000111000100    0100000111000101    0100000111000110    0100000111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16835 - 16839

  --0100000111001000    0100000111001001    0100000111001010    0100000111001011    0100000111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16840 - 16844

  --0100000111001101    0100000111001110    0100000111001111    0100000111010000    0100000111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16845 - 16849

  --0100000111010010    0100000111010011    0100000111010100    0100000111010101    0100000111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16850 - 16854

  --0100000111010111    0100000111011000    0100000111011001    0100000111011010    0100000111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16855 - 16859

  --0100000111011100    0100000111011101    0100000111011110    0100000111011111    0100000111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16860 - 16864

  --0100000111100001    0100000111100010    0100000111100011    0100000111100100    0100000111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16865 - 16869

  --0100000111100110    0100000111100111    0100000111101000    0100000111101001    0100000111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16870 - 16874

  --0100000111101011    0100000111101100    0100000111101101    0100000111101110    0100000111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16875 - 16879

  --0100000111110000    0100000111110001    0100000111110010    0100000111110011    0100000111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16880 - 16884

  --0100000111110101    0100000111110110    0100000111110111    0100000111111000    0100000111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16885 - 16889

  --0100000111111010    0100000111111011    0100000111111100    0100000111111101    0100000111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16890 - 16894

  --0100000111111111    0100001000000000    0100001000000001    0100001000000010    0100001000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16895 - 16899

  --0100001000000100    0100001000000101    0100001000000110    0100001000000111    0100001000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16900 - 16904

  --0100001000001001    0100001000001010    0100001000001011    0100001000001100    0100001000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16905 - 16909

  --0100001000001110    0100001000001111    0100001000010000    0100001000010001    0100001000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16910 - 16914

  --0100001000010011    0100001000010100    0100001000010101    0100001000010110    0100001000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16915 - 16919

  --0100001000011000    0100001000011001    0100001000011010    0100001000011011    0100001000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16920 - 16924

  --0100001000011101    0100001000011110    0100001000011111    0100001000100000    0100001000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16925 - 16929

  --0100001000100010    0100001000100011    0100001000100100    0100001000100101    0100001000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16930 - 16934

  --0100001000100111    0100001000101000    0100001000101001    0100001000101010    0100001000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16935 - 16939

  --0100001000101100    0100001000101101    0100001000101110    0100001000101111    0100001000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16940 - 16944

  --0100001000110001    0100001000110010    0100001000110011    0100001000110100    0100001000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16945 - 16949

  --0100001000110110    0100001000110111    0100001000111000    0100001000111001    0100001000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16950 - 16954

  --0100001000111011    0100001000111100    0100001000111101    0100001000111110    0100001000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16955 - 16959

  --0100001001000000    0100001001000001    0100001001000010    0100001001000011    0100001001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16960 - 16964

  --0100001001000101    0100001001000110    0100001001000111    0100001001001000    0100001001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16965 - 16969

  --0100001001001010    0100001001001011    0100001001001100    0100001001001101    0100001001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16970 - 16974

  --0100001001001111    0100001001010000    0100001001010001    0100001001010010    0100001001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16975 - 16979

  --0100001001010100    0100001001010101    0100001001010110    0100001001010111    0100001001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16980 - 16984

  --0100001001011001    0100001001011010    0100001001011011    0100001001011100    0100001001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16985 - 16989

  --0100001001011110    0100001001011111    0100001001100000    0100001001100001    0100001001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16990 - 16994

  --0100001001100011    0100001001100100    0100001001100101    0100001001100110    0100001001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 16995 - 16999

  --0100001001101000    0100001001101001    0100001001101010    0100001001101011    0100001001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17000 - 17004

  --0100001001101101    0100001001101110    0100001001101111    0100001001110000    0100001001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17005 - 17009

  --0100001001110010    0100001001110011    0100001001110100    0100001001110101    0100001001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17010 - 17014

  --0100001001110111    0100001001111000    0100001001111001    0100001001111010    0100001001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17015 - 17019

  --0100001001111100    0100001001111101    0100001001111110    0100001001111111    0100001010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17020 - 17024

  --0100001010000001    0100001010000010    0100001010000011    0100001010000100    0100001010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17025 - 17029

  --0100001010000110    0100001010000111    0100001010001000    0100001010001001    0100001010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17030 - 17034

  --0100001010001011    0100001010001100    0100001010001101    0100001010001110    0100001010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17035 - 17039

  --0100001010010000    0100001010010001    0100001010010010    0100001010010011    0100001010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17040 - 17044

  --0100001010010101    0100001010010110    0100001010010111    0100001010011000    0100001010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17045 - 17049

  --0100001010011010    0100001010011011    0100001010011100    0100001010011101    0100001010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17050 - 17054

  --0100001010011111    0100001010100000    0100001010100001    0100001010100010    0100001010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17055 - 17059

  --0100001010100100    0100001010100101    0100001010100110    0100001010100111    0100001010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17060 - 17064

  --0100001010101001    0100001010101010    0100001010101011    0100001010101100    0100001010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17065 - 17069

  --0100001010101110    0100001010101111    0100001010110000    0100001010110001    0100001010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17070 - 17074

  --0100001010110011    0100001010110100    0100001010110101    0100001010110110    0100001010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17075 - 17079

  --0100001010111000    0100001010111001    0100001010111010    0100001010111011    0100001010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17080 - 17084

  --0100001010111101    0100001010111110    0100001010111111    0100001011000000    0100001011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17085 - 17089

  --0100001011000010    0100001011000011    0100001011000100    0100001011000101    0100001011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17090 - 17094

  --0100001011000111    0100001011001000    0100001011001001    0100001011001010    0100001011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17095 - 17099

  --0100001011001100    0100001011001101    0100001011001110    0100001011001111    0100001011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17100 - 17104

  --0100001011010001    0100001011010010    0100001011010011    0100001011010100    0100001011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17105 - 17109

  --0100001011010110    0100001011010111    0100001011011000    0100001011011001    0100001011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17110 - 17114

  --0100001011011011    0100001011011100    0100001011011101    0100001011011110    0100001011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17115 - 17119

  --0100001011100000    0100001011100001    0100001011100010    0100001011100011    0100001011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17120 - 17124

  --0100001011100101    0100001011100110    0100001011100111    0100001011101000    0100001011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17125 - 17129

  --0100001011101010    0100001011101011    0100001011101100    0100001011101101    0100001011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17130 - 17134

  --0100001011101111    0100001011110000    0100001011110001    0100001011110010    0100001011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17135 - 17139

  --0100001011110100    0100001011110101    0100001011110110    0100001011110111    0100001011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17140 - 17144

  --0100001011111001    0100001011111010    0100001011111011    0100001011111100    0100001011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17145 - 17149

  --0100001011111110    0100001011111111    0100001100000000    0100001100000001    0100001100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17150 - 17154

  --0100001100000011    0100001100000100    0100001100000101    0100001100000110    0100001100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17155 - 17159

  --0100001100001000    0100001100001001    0100001100001010    0100001100001011    0100001100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17160 - 17164

  --0100001100001101    0100001100001110    0100001100001111    0100001100010000    0100001100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17165 - 17169

  --0100001100010010    0100001100010011    0100001100010100    0100001100010101    0100001100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17170 - 17174

  --0100001100010111    0100001100011000    0100001100011001    0100001100011010    0100001100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17175 - 17179

  --0100001100011100    0100001100011101    0100001100011110    0100001100011111    0100001100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17180 - 17184

  --0100001100100001    0100001100100010    0100001100100011    0100001100100100    0100001100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17185 - 17189

  --0100001100100110    0100001100100111    0100001100101000    0100001100101001    0100001100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17190 - 17194

  --0100001100101011    0100001100101100    0100001100101101    0100001100101110    0100001100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17195 - 17199

  --0100001100110000    0100001100110001    0100001100110010    0100001100110011    0100001100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17200 - 17204

  --0100001100110101    0100001100110110    0100001100110111    0100001100111000    0100001100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17205 - 17209

  --0100001100111010    0100001100111011    0100001100111100    0100001100111101    0100001100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17210 - 17214

  --0100001100111111    0100001101000000    0100001101000001    0100001101000010    0100001101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17215 - 17219

  --0100001101000100    0100001101000101    0100001101000110    0100001101000111    0100001101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17220 - 17224

  --0100001101001001    0100001101001010    0100001101001011    0100001101001100    0100001101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17225 - 17229

  --0100001101001110    0100001101001111    0100001101010000    0100001101010001    0100001101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17230 - 17234

  --0100001101010011    0100001101010100    0100001101010101    0100001101010110    0100001101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17235 - 17239

  --0100001101011000    0100001101011001    0100001101011010    0100001101011011    0100001101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17240 - 17244

  --0100001101011101    0100001101011110    0100001101011111    0100001101100000    0100001101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17245 - 17249

  --0100001101100010    0100001101100011    0100001101100100    0100001101100101    0100001101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17250 - 17254

  --0100001101100111    0100001101101000    0100001101101001    0100001101101010    0100001101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17255 - 17259

  --0100001101101100    0100001101101101    0100001101101110    0100001101101111    0100001101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17260 - 17264

  --0100001101110001    0100001101110010    0100001101110011    0100001101110100    0100001101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17265 - 17269

  --0100001101110110    0100001101110111    0100001101111000    0100001101111001    0100001101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17270 - 17274

  --0100001101111011    0100001101111100    0100001101111101    0100001101111110    0100001101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17275 - 17279

  --0100001110000000    0100001110000001    0100001110000010    0100001110000011    0100001110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17280 - 17284

  --0100001110000101    0100001110000110    0100001110000111    0100001110001000    0100001110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17285 - 17289

  --0100001110001010    0100001110001011    0100001110001100    0100001110001101    0100001110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17290 - 17294

  --0100001110001111    0100001110010000    0100001110010001    0100001110010010    0100001110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17295 - 17299

  --0100001110010100    0100001110010101    0100001110010110    0100001110010111    0100001110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17300 - 17304

  --0100001110011001    0100001110011010    0100001110011011    0100001110011100    0100001110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17305 - 17309

  --0100001110011110    0100001110011111    0100001110100000    0100001110100001    0100001110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17310 - 17314

  --0100001110100011    0100001110100100    0100001110100101    0100001110100110    0100001110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17315 - 17319

  --0100001110101000    0100001110101001    0100001110101010    0100001110101011    0100001110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17320 - 17324

  --0100001110101101    0100001110101110    0100001110101111    0100001110110000    0100001110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17325 - 17329

  --0100001110110010    0100001110110011    0100001110110100    0100001110110101    0100001110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17330 - 17334

  --0100001110110111    0100001110111000    0100001110111001    0100001110111010    0100001110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17335 - 17339

  --0100001110111100    0100001110111101    0100001110111110    0100001110111111    0100001111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17340 - 17344

  --0100001111000001    0100001111000010    0100001111000011    0100001111000100    0100001111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17345 - 17349

  --0100001111000110    0100001111000111    0100001111001000    0100001111001001    0100001111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17350 - 17354

  --0100001111001011    0100001111001100    0100001111001101    0100001111001110    0100001111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17355 - 17359

  --0100001111010000    0100001111010001    0100001111010010    0100001111010011    0100001111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17360 - 17364

  --0100001111010101    0100001111010110    0100001111010111    0100001111011000    0100001111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17365 - 17369

  --0100001111011010    0100001111011011    0100001111011100    0100001111011101    0100001111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17370 - 17374

  --0100001111011111    0100001111100000    0100001111100001    0100001111100010    0100001111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17375 - 17379

  --0100001111100100    0100001111100101    0100001111100110    0100001111100111    0100001111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17380 - 17384

  --0100001111101001    0100001111101010    0100001111101011    0100001111101100    0100001111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17385 - 17389

  --0100001111101110    0100001111101111    0100001111110000    0100001111110001    0100001111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17390 - 17394

  --0100001111110011    0100001111110100    0100001111110101    0100001111110110    0100001111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17395 - 17399

  --0100001111111000    0100001111111001    0100001111111010    0100001111111011    0100001111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17400 - 17404

  --0100001111111101    0100001111111110    0100001111111111    0100010000000000    0100010000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17405 - 17409

  --0100010000000010    0100010000000011    0100010000000100    0100010000000101    0100010000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17410 - 17414

  --0100010000000111    0100010000001000    0100010000001001    0100010000001010    0100010000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17415 - 17419

  --0100010000001100    0100010000001101    0100010000001110    0100010000001111    0100010000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17420 - 17424

  --0100010000010001    0100010000010010    0100010000010011    0100010000010100    0100010000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17425 - 17429

  --0100010000010110    0100010000010111    0100010000011000    0100010000011001    0100010000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17430 - 17434

  --0100010000011011    0100010000011100    0100010000011101    0100010000011110    0100010000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17435 - 17439

  --0100010000100000    0100010000100001    0100010000100010    0100010000100011    0100010000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17440 - 17444

  --0100010000100101    0100010000100110    0100010000100111    0100010000101000    0100010000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17445 - 17449

  --0100010000101010    0100010000101011    0100010000101100    0100010000101101    0100010000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17450 - 17454

  --0100010000101111    0100010000110000    0100010000110001    0100010000110010    0100010000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17455 - 17459

  --0100010000110100    0100010000110101    0100010000110110    0100010000110111    0100010000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17460 - 17464

  --0100010000111001    0100010000111010    0100010000111011    0100010000111100    0100010000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17465 - 17469

  --0100010000111110    0100010000111111    0100010001000000    0100010001000001    0100010001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17470 - 17474

  --0100010001000011    0100010001000100    0100010001000101    0100010001000110    0100010001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17475 - 17479

  --0100010001001000    0100010001001001    0100010001001010    0100010001001011    0100010001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17480 - 17484

  --0100010001001101    0100010001001110    0100010001001111    0100010001010000    0100010001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17485 - 17489

  --0100010001010010    0100010001010011    0100010001010100    0100010001010101    0100010001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17490 - 17494

  --0100010001010111    0100010001011000    0100010001011001    0100010001011010    0100010001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17495 - 17499

  --0100010001011100    0100010001011101    0100010001011110    0100010001011111    0100010001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17500 - 17504

  --0100010001100001    0100010001100010    0100010001100011    0100010001100100    0100010001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17505 - 17509

  --0100010001100110    0100010001100111    0100010001101000    0100010001101001    0100010001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17510 - 17514

  --0100010001101011    0100010001101100    0100010001101101    0100010001101110    0100010001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17515 - 17519

  --0100010001110000    0100010001110001    0100010001110010    0100010001110011    0100010001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17520 - 17524

  --0100010001110101    0100010001110110    0100010001110111    0100010001111000    0100010001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17525 - 17529

  --0100010001111010    0100010001111011    0100010001111100    0100010001111101    0100010001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17530 - 17534

  --0100010001111111    0100010010000000    0100010010000001    0100010010000010    0100010010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17535 - 17539

  --0100010010000100    0100010010000101    0100010010000110    0100010010000111    0100010010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17540 - 17544

  --0100010010001001    0100010010001010    0100010010001011    0100010010001100    0100010010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17545 - 17549

  --0100010010001110    0100010010001111    0100010010010000    0100010010010001    0100010010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17550 - 17554

  --0100010010010011    0100010010010100    0100010010010101    0100010010010110    0100010010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17555 - 17559

  --0100010010011000    0100010010011001    0100010010011010    0100010010011011    0100010010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17560 - 17564

  --0100010010011101    0100010010011110    0100010010011111    0100010010100000    0100010010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17565 - 17569

  --0100010010100010    0100010010100011    0100010010100100    0100010010100101    0100010010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17570 - 17574

  --0100010010100111    0100010010101000    0100010010101001    0100010010101010    0100010010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17575 - 17579

  --0100010010101100    0100010010101101    0100010010101110    0100010010101111    0100010010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17580 - 17584

  --0100010010110001    0100010010110010    0100010010110011    0100010010110100    0100010010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17585 - 17589

  --0100010010110110    0100010010110111    0100010010111000    0100010010111001    0100010010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17590 - 17594

  --0100010010111011    0100010010111100    0100010010111101    0100010010111110    0100010010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17595 - 17599

  --0100010011000000    0100010011000001    0100010011000010    0100010011000011    0100010011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17600 - 17604

  --0100010011000101    0100010011000110    0100010011000111    0100010011001000    0100010011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17605 - 17609

  --0100010011001010    0100010011001011    0100010011001100    0100010011001101    0100010011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17610 - 17614

  --0100010011001111    0100010011010000    0100010011010001    0100010011010010    0100010011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17615 - 17619

  --0100010011010100    0100010011010101    0100010011010110    0100010011010111    0100010011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17620 - 17624

  --0100010011011001    0100010011011010    0100010011011011    0100010011011100    0100010011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17625 - 17629

  --0100010011011110    0100010011011111    0100010011100000    0100010011100001    0100010011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17630 - 17634

  --0100010011100011    0100010011100100    0100010011100101    0100010011100110    0100010011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17635 - 17639

  --0100010011101000    0100010011101001    0100010011101010    0100010011101011    0100010011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17640 - 17644

  --0100010011101101    0100010011101110    0100010011101111    0100010011110000    0100010011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17645 - 17649

  --0100010011110010    0100010011110011    0100010011110100    0100010011110101    0100010011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17650 - 17654

  --0100010011110111    0100010011111000    0100010011111001    0100010011111010    0100010011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17655 - 17659

  --0100010011111100    0100010011111101    0100010011111110    0100010011111111    0100010100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17660 - 17664

  --0100010100000001    0100010100000010    0100010100000011    0100010100000100    0100010100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17665 - 17669

  --0100010100000110    0100010100000111    0100010100001000    0100010100001001    0100010100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17670 - 17674

  --0100010100001011    0100010100001100    0100010100001101    0100010100001110    0100010100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17675 - 17679

  --0100010100010000    0100010100010001    0100010100010010    0100010100010011    0100010100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17680 - 17684

  --0100010100010101    0100010100010110    0100010100010111    0100010100011000    0100010100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17685 - 17689

  --0100010100011010    0100010100011011    0100010100011100    0100010100011101    0100010100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17690 - 17694

  --0100010100011111    0100010100100000    0100010100100001    0100010100100010    0100010100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17695 - 17699

  --0100010100100100    0100010100100101    0100010100100110    0100010100100111    0100010100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17700 - 17704

  --0100010100101001    0100010100101010    0100010100101011    0100010100101100    0100010100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17705 - 17709

  --0100010100101110    0100010100101111    0100010100110000    0100010100110001    0100010100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17710 - 17714

  --0100010100110011    0100010100110100    0100010100110101    0100010100110110    0100010100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17715 - 17719

  --0100010100111000    0100010100111001    0100010100111010    0100010100111011    0100010100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17720 - 17724

  --0100010100111101    0100010100111110    0100010100111111    0100010101000000    0100010101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17725 - 17729

  --0100010101000010    0100010101000011    0100010101000100    0100010101000101    0100010101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17730 - 17734

  --0100010101000111    0100010101001000    0100010101001001    0100010101001010    0100010101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17735 - 17739

  --0100010101001100    0100010101001101    0100010101001110    0100010101001111    0100010101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17740 - 17744

  --0100010101010001    0100010101010010    0100010101010011    0100010101010100    0100010101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17745 - 17749

  --0100010101010110    0100010101010111    0100010101011000    0100010101011001    0100010101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17750 - 17754

  --0100010101011011    0100010101011100    0100010101011101    0100010101011110    0100010101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17755 - 17759

  --0100010101100000    0100010101100001    0100010101100010    0100010101100011    0100010101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17760 - 17764

  --0100010101100101    0100010101100110    0100010101100111    0100010101101000    0100010101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17765 - 17769

  --0100010101101010    0100010101101011    0100010101101100    0100010101101101    0100010101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17770 - 17774

  --0100010101101111    0100010101110000    0100010101110001    0100010101110010    0100010101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17775 - 17779

  --0100010101110100    0100010101110101    0100010101110110    0100010101110111    0100010101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17780 - 17784

  --0100010101111001    0100010101111010    0100010101111011    0100010101111100    0100010101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17785 - 17789

  --0100010101111110    0100010101111111    0100010110000000    0100010110000001    0100010110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17790 - 17794

  --0100010110000011    0100010110000100    0100010110000101    0100010110000110    0100010110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17795 - 17799

  --0100010110001000    0100010110001001    0100010110001010    0100010110001011    0100010110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17800 - 17804

  --0100010110001101    0100010110001110    0100010110001111    0100010110010000    0100010110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17805 - 17809

  --0100010110010010    0100010110010011    0100010110010100    0100010110010101    0100010110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17810 - 17814

  --0100010110010111    0100010110011000    0100010110011001    0100010110011010    0100010110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17815 - 17819

  --0100010110011100    0100010110011101    0100010110011110    0100010110011111    0100010110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17820 - 17824

  --0100010110100001    0100010110100010    0100010110100011    0100010110100100    0100010110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17825 - 17829

  --0100010110100110    0100010110100111    0100010110101000    0100010110101001    0100010110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17830 - 17834

  --0100010110101011    0100010110101100    0100010110101101    0100010110101110    0100010110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17835 - 17839

  --0100010110110000    0100010110110001    0100010110110010    0100010110110011    0100010110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17840 - 17844

  --0100010110110101    0100010110110110    0100010110110111    0100010110111000    0100010110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17845 - 17849

  --0100010110111010    0100010110111011    0100010110111100    0100010110111101    0100010110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17850 - 17854

  --0100010110111111    0100010111000000    0100010111000001    0100010111000010    0100010111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17855 - 17859

  --0100010111000100    0100010111000101    0100010111000110    0100010111000111    0100010111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17860 - 17864

  --0100010111001001    0100010111001010    0100010111001011    0100010111001100    0100010111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17865 - 17869

  --0100010111001110    0100010111001111    0100010111010000    0100010111010001    0100010111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17870 - 17874

  --0100010111010011    0100010111010100    0100010111010101    0100010111010110    0100010111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17875 - 17879

  --0100010111011000    0100010111011001    0100010111011010    0100010111011011    0100010111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17880 - 17884

  --0100010111011101    0100010111011110    0100010111011111    0100010111100000    0100010111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17885 - 17889

  --0100010111100010    0100010111100011    0100010111100100    0100010111100101    0100010111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17890 - 17894

  --0100010111100111    0100010111101000    0100010111101001    0100010111101010    0100010111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17895 - 17899

  --0100010111101100    0100010111101101    0100010111101110    0100010111101111    0100010111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17900 - 17904

  --0100010111110001    0100010111110010    0100010111110011    0100010111110100    0100010111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17905 - 17909

  --0100010111110110    0100010111110111    0100010111111000    0100010111111001    0100010111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17910 - 17914

  --0100010111111011    0100010111111100    0100010111111101    0100010111111110    0100010111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17915 - 17919

  --0100011000000000    0100011000000001    0100011000000010    0100011000000011    0100011000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17920 - 17924

  --0100011000000101    0100011000000110    0100011000000111    0100011000001000    0100011000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17925 - 17929

  --0100011000001010    0100011000001011    0100011000001100    0100011000001101    0100011000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17930 - 17934

  --0100011000001111    0100011000010000    0100011000010001    0100011000010010    0100011000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17935 - 17939

  --0100011000010100    0100011000010101    0100011000010110    0100011000010111    0100011000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17940 - 17944

  --0100011000011001    0100011000011010    0100011000011011    0100011000011100    0100011000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17945 - 17949

  --0100011000011110    0100011000011111    0100011000100000    0100011000100001    0100011000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17950 - 17954

  --0100011000100011    0100011000100100    0100011000100101    0100011000100110    0100011000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17955 - 17959

  --0100011000101000    0100011000101001    0100011000101010    0100011000101011    0100011000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17960 - 17964

  --0100011000101101    0100011000101110    0100011000101111    0100011000110000    0100011000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17965 - 17969

  --0100011000110010    0100011000110011    0100011000110100    0100011000110101    0100011000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17970 - 17974

  --0100011000110111    0100011000111000    0100011000111001    0100011000111010    0100011000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17975 - 17979

  --0100011000111100    0100011000111101    0100011000111110    0100011000111111    0100011001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17980 - 17984

  --0100011001000001    0100011001000010    0100011001000011    0100011001000100    0100011001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17985 - 17989

  --0100011001000110    0100011001000111    0100011001001000    0100011001001001    0100011001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17990 - 17994

  --0100011001001011    0100011001001100    0100011001001101    0100011001001110    0100011001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 17995 - 17999

  --0100011001010000    0100011001010001    0100011001010010    0100011001010011    0100011001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18000 - 18004

  --0100011001010101    0100011001010110    0100011001010111    0100011001011000    0100011001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18005 - 18009

  --0100011001011010    0100011001011011    0100011001011100    0100011001011101    0100011001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18010 - 18014

  --0100011001011111    0100011001100000    0100011001100001    0100011001100010    0100011001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18015 - 18019

  --0100011001100100    0100011001100101    0100011001100110    0100011001100111    0100011001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18020 - 18024

  --0100011001101001    0100011001101010    0100011001101011    0100011001101100    0100011001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18025 - 18029

  --0100011001101110    0100011001101111    0100011001110000    0100011001110001    0100011001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18030 - 18034

  --0100011001110011    0100011001110100    0100011001110101    0100011001110110    0100011001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18035 - 18039

  --0100011001111000    0100011001111001    0100011001111010    0100011001111011    0100011001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18040 - 18044

  --0100011001111101    0100011001111110    0100011001111111    0100011010000000    0100011010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18045 - 18049

  --0100011010000010    0100011010000011    0100011010000100    0100011010000101    0100011010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18050 - 18054

  --0100011010000111    0100011010001000    0100011010001001    0100011010001010    0100011010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18055 - 18059

  --0100011010001100    0100011010001101    0100011010001110    0100011010001111    0100011010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18060 - 18064

  --0100011010010001    0100011010010010    0100011010010011    0100011010010100    0100011010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18065 - 18069

  --0100011010010110    0100011010010111    0100011010011000    0100011010011001    0100011010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18070 - 18074

  --0100011010011011    0100011010011100    0100011010011101    0100011010011110    0100011010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18075 - 18079

  --0100011010100000    0100011010100001    0100011010100010    0100011010100011    0100011010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18080 - 18084

  --0100011010100101    0100011010100110    0100011010100111    0100011010101000    0100011010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18085 - 18089

  --0100011010101010    0100011010101011    0100011010101100    0100011010101101    0100011010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18090 - 18094

  --0100011010101111    0100011010110000    0100011010110001    0100011010110010    0100011010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18095 - 18099

  --0100011010110100    0100011010110101    0100011010110110    0100011010110111    0100011010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18100 - 18104

  --0100011010111001    0100011010111010    0100011010111011    0100011010111100    0100011010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18105 - 18109

  --0100011010111110    0100011010111111    0100011011000000    0100011011000001    0100011011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18110 - 18114

  --0100011011000011    0100011011000100    0100011011000101    0100011011000110    0100011011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18115 - 18119

  --0100011011001000    0100011011001001    0100011011001010    0100011011001011    0100011011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18120 - 18124

  --0100011011001101    0100011011001110    0100011011001111    0100011011010000    0100011011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18125 - 18129

  --0100011011010010    0100011011010011    0100011011010100    0100011011010101    0100011011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18130 - 18134

  --0100011011010111    0100011011011000    0100011011011001    0100011011011010    0100011011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18135 - 18139

  --0100011011011100    0100011011011101    0100011011011110    0100011011011111    0100011011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18140 - 18144

  --0100011011100001    0100011011100010    0100011011100011    0100011011100100    0100011011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18145 - 18149

  --0100011011100110    0100011011100111    0100011011101000    0100011011101001    0100011011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18150 - 18154

  --0100011011101011    0100011011101100    0100011011101101    0100011011101110    0100011011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18155 - 18159

  --0100011011110000    0100011011110001    0100011011110010    0100011011110011    0100011011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18160 - 18164

  --0100011011110101    0100011011110110    0100011011110111    0100011011111000    0100011011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18165 - 18169

  --0100011011111010    0100011011111011    0100011011111100    0100011011111101    0100011011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18170 - 18174

  --0100011011111111    0100011100000000    0100011100000001    0100011100000010    0100011100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18175 - 18179

  --0100011100000100    0100011100000101    0100011100000110    0100011100000111    0100011100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18180 - 18184

  --0100011100001001    0100011100001010    0100011100001011    0100011100001100    0100011100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18185 - 18189

  --0100011100001110    0100011100001111    0100011100010000    0100011100010001    0100011100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18190 - 18194

  --0100011100010011    0100011100010100    0100011100010101    0100011100010110    0100011100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18195 - 18199

  --0100011100011000    0100011100011001    0100011100011010    0100011100011011    0100011100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18200 - 18204

  --0100011100011101    0100011100011110    0100011100011111    0100011100100000    0100011100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18205 - 18209

  --0100011100100010    0100011100100011    0100011100100100    0100011100100101    0100011100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18210 - 18214

  --0100011100100111    0100011100101000    0100011100101001    0100011100101010    0100011100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18215 - 18219

  --0100011100101100    0100011100101101    0100011100101110    0100011100101111    0100011100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18220 - 18224

  --0100011100110001    0100011100110010    0100011100110011    0100011100110100    0100011100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18225 - 18229

  --0100011100110110    0100011100110111    0100011100111000    0100011100111001    0100011100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18230 - 18234

  --0100011100111011    0100011100111100    0100011100111101    0100011100111110    0100011100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18235 - 18239

  --0100011101000000    0100011101000001    0100011101000010    0100011101000011    0100011101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18240 - 18244

  --0100011101000101    0100011101000110    0100011101000111    0100011101001000    0100011101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18245 - 18249

  --0100011101001010    0100011101001011    0100011101001100    0100011101001101    0100011101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18250 - 18254

  --0100011101001111    0100011101010000    0100011101010001    0100011101010010    0100011101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18255 - 18259

  --0100011101010100    0100011101010101    0100011101010110    0100011101010111    0100011101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18260 - 18264

  --0100011101011001    0100011101011010    0100011101011011    0100011101011100    0100011101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18265 - 18269

  --0100011101011110    0100011101011111    0100011101100000    0100011101100001    0100011101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18270 - 18274

  --0100011101100011    0100011101100100    0100011101100101    0100011101100110    0100011101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18275 - 18279

  --0100011101101000    0100011101101001    0100011101101010    0100011101101011    0100011101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18280 - 18284

  --0100011101101101    0100011101101110    0100011101101111    0100011101110000    0100011101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18285 - 18289

  --0100011101110010    0100011101110011    0100011101110100    0100011101110101    0100011101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18290 - 18294

  --0100011101110111    0100011101111000    0100011101111001    0100011101111010    0100011101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18295 - 18299

  --0100011101111100    0100011101111101    0100011101111110    0100011101111111    0100011110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18300 - 18304

  --0100011110000001    0100011110000010    0100011110000011    0100011110000100    0100011110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18305 - 18309

  --0100011110000110    0100011110000111    0100011110001000    0100011110001001    0100011110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18310 - 18314

  --0100011110001011    0100011110001100    0100011110001101    0100011110001110    0100011110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18315 - 18319

  --0100011110010000    0100011110010001    0100011110010010    0100011110010011    0100011110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18320 - 18324

  --0100011110010101    0100011110010110    0100011110010111    0100011110011000    0100011110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18325 - 18329

  --0100011110011010    0100011110011011    0100011110011100    0100011110011101    0100011110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18330 - 18334

  --0100011110011111    0100011110100000    0100011110100001    0100011110100010    0100011110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18335 - 18339

  --0100011110100100    0100011110100101    0100011110100110    0100011110100111    0100011110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18340 - 18344

  --0100011110101001    0100011110101010    0100011110101011    0100011110101100    0100011110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18345 - 18349

  --0100011110101110    0100011110101111    0100011110110000    0100011110110001    0100011110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18350 - 18354

  --0100011110110011    0100011110110100    0100011110110101    0100011110110110    0100011110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18355 - 18359

  --0100011110111000    0100011110111001    0100011110111010    0100011110111011    0100011110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18360 - 18364

  --0100011110111101    0100011110111110    0100011110111111    0100011111000000    0100011111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18365 - 18369

  --0100011111000010    0100011111000011    0100011111000100    0100011111000101    0100011111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18370 - 18374

  --0100011111000111    0100011111001000    0100011111001001    0100011111001010    0100011111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18375 - 18379

  --0100011111001100    0100011111001101    0100011111001110    0100011111001111    0100011111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18380 - 18384

  --0100011111010001    0100011111010010    0100011111010011    0100011111010100    0100011111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18385 - 18389

  --0100011111010110    0100011111010111    0100011111011000    0100011111011001    0100011111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18390 - 18394

  --0100011111011011    0100011111011100    0100011111011101    0100011111011110    0100011111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18395 - 18399

  --0100011111100000    0100011111100001    0100011111100010    0100011111100011    0100011111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18400 - 18404

  --0100011111100101    0100011111100110    0100011111100111    0100011111101000    0100011111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18405 - 18409

  --0100011111101010    0100011111101011    0100011111101100    0100011111101101    0100011111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18410 - 18414

  --0100011111101111    0100011111110000    0100011111110001    0100011111110010    0100011111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18415 - 18419

  --0100011111110100    0100011111110101    0100011111110110    0100011111110111    0100011111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18420 - 18424

  --0100011111111001    0100011111111010    0100011111111011    0100011111111100    0100011111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18425 - 18429

  --0100011111111110    0100011111111111    0100100000000000    0100100000000001    0100100000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18430 - 18434

  --0100100000000011    0100100000000100    0100100000000101    0100100000000110    0100100000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18435 - 18439

  --0100100000001000    0100100000001001    0100100000001010    0100100000001011    0100100000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18440 - 18444

  --0100100000001101    0100100000001110    0100100000001111    0100100000010000    0100100000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18445 - 18449

  --0100100000010010    0100100000010011    0100100000010100    0100100000010101    0100100000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18450 - 18454

  --0100100000010111    0100100000011000    0100100000011001    0100100000011010    0100100000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18455 - 18459

  --0100100000011100    0100100000011101    0100100000011110    0100100000011111    0100100000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18460 - 18464

  --0100100000100001    0100100000100010    0100100000100011    0100100000100100    0100100000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18465 - 18469

  --0100100000100110    0100100000100111    0100100000101000    0100100000101001    0100100000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18470 - 18474

  --0100100000101011    0100100000101100    0100100000101101    0100100000101110    0100100000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18475 - 18479

  --0100100000110000    0100100000110001    0100100000110010    0100100000110011    0100100000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18480 - 18484

  --0100100000110101    0100100000110110    0100100000110111    0100100000111000    0100100000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18485 - 18489

  --0100100000111010    0100100000111011    0100100000111100    0100100000111101    0100100000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18490 - 18494

  --0100100000111111    0100100001000000    0100100001000001    0100100001000010    0100100001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18495 - 18499

  --0100100001000100    0100100001000101    0100100001000110    0100100001000111    0100100001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18500 - 18504

  --0100100001001001    0100100001001010    0100100001001011    0100100001001100    0100100001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18505 - 18509

  --0100100001001110    0100100001001111    0100100001010000    0100100001010001    0100100001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18510 - 18514

  --0100100001010011    0100100001010100    0100100001010101    0100100001010110    0100100001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18515 - 18519

  --0100100001011000    0100100001011001    0100100001011010    0100100001011011    0100100001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18520 - 18524

  --0100100001011101    0100100001011110    0100100001011111    0100100001100000    0100100001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18525 - 18529

  --0100100001100010    0100100001100011    0100100001100100    0100100001100101    0100100001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18530 - 18534

  --0100100001100111    0100100001101000    0100100001101001    0100100001101010    0100100001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18535 - 18539

  --0100100001101100    0100100001101101    0100100001101110    0100100001101111    0100100001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18540 - 18544

  --0100100001110001    0100100001110010    0100100001110011    0100100001110100    0100100001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18545 - 18549

  --0100100001110110    0100100001110111    0100100001111000    0100100001111001    0100100001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18550 - 18554

  --0100100001111011    0100100001111100    0100100001111101    0100100001111110    0100100001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18555 - 18559

  --0100100010000000    0100100010000001    0100100010000010    0100100010000011    0100100010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18560 - 18564

  --0100100010000101    0100100010000110    0100100010000111    0100100010001000    0100100010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18565 - 18569

  --0100100010001010    0100100010001011    0100100010001100    0100100010001101    0100100010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18570 - 18574

  --0100100010001111    0100100010010000    0100100010010001    0100100010010010    0100100010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18575 - 18579

  --0100100010010100    0100100010010101    0100100010010110    0100100010010111    0100100010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18580 - 18584

  --0100100010011001    0100100010011010    0100100010011011    0100100010011100    0100100010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18585 - 18589

  --0100100010011110    0100100010011111    0100100010100000    0100100010100001    0100100010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18590 - 18594

  --0100100010100011    0100100010100100    0100100010100101    0100100010100110    0100100010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18595 - 18599

  --0100100010101000    0100100010101001    0100100010101010    0100100010101011    0100100010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18600 - 18604

  --0100100010101101    0100100010101110    0100100010101111    0100100010110000    0100100010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18605 - 18609

  --0100100010110010    0100100010110011    0100100010110100    0100100010110101    0100100010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18610 - 18614

  --0100100010110111    0100100010111000    0100100010111001    0100100010111010    0100100010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18615 - 18619

  --0100100010111100    0100100010111101    0100100010111110    0100100010111111    0100100011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18620 - 18624

  --0100100011000001    0100100011000010    0100100011000011    0100100011000100    0100100011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18625 - 18629

  --0100100011000110    0100100011000111    0100100011001000    0100100011001001    0100100011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18630 - 18634

  --0100100011001011    0100100011001100    0100100011001101    0100100011001110    0100100011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18635 - 18639

  --0100100011010000    0100100011010001    0100100011010010    0100100011010011    0100100011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18640 - 18644

  --0100100011010101    0100100011010110    0100100011010111    0100100011011000    0100100011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18645 - 18649

  --0100100011011010    0100100011011011    0100100011011100    0100100011011101    0100100011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18650 - 18654

  --0100100011011111    0100100011100000    0100100011100001    0100100011100010    0100100011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18655 - 18659

  --0100100011100100    0100100011100101    0100100011100110    0100100011100111    0100100011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18660 - 18664

  --0100100011101001    0100100011101010    0100100011101011    0100100011101100    0100100011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18665 - 18669

  --0100100011101110    0100100011101111    0100100011110000    0100100011110001    0100100011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18670 - 18674

  --0100100011110011    0100100011110100    0100100011110101    0100100011110110    0100100011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18675 - 18679

  --0100100011111000    0100100011111001    0100100011111010    0100100011111011    0100100011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18680 - 18684

  --0100100011111101    0100100011111110    0100100011111111    0100100100000000    0100100100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18685 - 18689

  --0100100100000010    0100100100000011    0100100100000100    0100100100000101    0100100100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18690 - 18694

  --0100100100000111    0100100100001000    0100100100001001    0100100100001010    0100100100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18695 - 18699

  --0100100100001100    0100100100001101    0100100100001110    0100100100001111    0100100100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18700 - 18704

  --0100100100010001    0100100100010010    0100100100010011    0100100100010100    0100100100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18705 - 18709

  --0100100100010110    0100100100010111    0100100100011000    0100100100011001    0100100100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18710 - 18714

  --0100100100011011    0100100100011100    0100100100011101    0100100100011110    0100100100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18715 - 18719

  --0100100100100000    0100100100100001    0100100100100010    0100100100100011    0100100100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18720 - 18724

  --0100100100100101    0100100100100110    0100100100100111    0100100100101000    0100100100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18725 - 18729

  --0100100100101010    0100100100101011    0100100100101100    0100100100101101    0100100100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18730 - 18734

  --0100100100101111    0100100100110000    0100100100110001    0100100100110010    0100100100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18735 - 18739

  --0100100100110100    0100100100110101    0100100100110110    0100100100110111    0100100100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18740 - 18744

  --0100100100111001    0100100100111010    0100100100111011    0100100100111100    0100100100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18745 - 18749

  --0100100100111110    0100100100111111    0100100101000000    0100100101000001    0100100101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18750 - 18754

  --0100100101000011    0100100101000100    0100100101000101    0100100101000110    0100100101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18755 - 18759

  --0100100101001000    0100100101001001    0100100101001010    0100100101001011    0100100101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18760 - 18764

  --0100100101001101    0100100101001110    0100100101001111    0100100101010000    0100100101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18765 - 18769

  --0100100101010010    0100100101010011    0100100101010100    0100100101010101    0100100101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18770 - 18774

  --0100100101010111    0100100101011000    0100100101011001    0100100101011010    0100100101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18775 - 18779

  --0100100101011100    0100100101011101    0100100101011110    0100100101011111    0100100101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18780 - 18784

  --0100100101100001    0100100101100010    0100100101100011    0100100101100100    0100100101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18785 - 18789

  --0100100101100110    0100100101100111    0100100101101000    0100100101101001    0100100101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18790 - 18794

  --0100100101101011    0100100101101100    0100100101101101    0100100101101110    0100100101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18795 - 18799

  --0100100101110000    0100100101110001    0100100101110010    0100100101110011    0100100101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18800 - 18804

  --0100100101110101    0100100101110110    0100100101110111    0100100101111000    0100100101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18805 - 18809

  --0100100101111010    0100100101111011    0100100101111100    0100100101111101    0100100101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18810 - 18814

  --0100100101111111    0100100110000000    0100100110000001    0100100110000010    0100100110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18815 - 18819

  --0100100110000100    0100100110000101    0100100110000110    0100100110000111    0100100110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18820 - 18824

  --0100100110001001    0100100110001010    0100100110001011    0100100110001100    0100100110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18825 - 18829

  --0100100110001110    0100100110001111    0100100110010000    0100100110010001    0100100110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18830 - 18834

  --0100100110010011    0100100110010100    0100100110010101    0100100110010110    0100100110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18835 - 18839

  --0100100110011000    0100100110011001    0100100110011010    0100100110011011    0100100110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18840 - 18844

  --0100100110011101    0100100110011110    0100100110011111    0100100110100000    0100100110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18845 - 18849

  --0100100110100010    0100100110100011    0100100110100100    0100100110100101    0100100110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18850 - 18854

  --0100100110100111    0100100110101000    0100100110101001    0100100110101010    0100100110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18855 - 18859

  --0100100110101100    0100100110101101    0100100110101110    0100100110101111    0100100110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18860 - 18864

  --0100100110110001    0100100110110010    0100100110110011    0100100110110100    0100100110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18865 - 18869

  --0100100110110110    0100100110110111    0100100110111000    0100100110111001    0100100110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18870 - 18874

  --0100100110111011    0100100110111100    0100100110111101    0100100110111110    0100100110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18875 - 18879

  --0100100111000000    0100100111000001    0100100111000010    0100100111000011    0100100111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18880 - 18884

  --0100100111000101    0100100111000110    0100100111000111    0100100111001000    0100100111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18885 - 18889

  --0100100111001010    0100100111001011    0100100111001100    0100100111001101    0100100111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18890 - 18894

  --0100100111001111    0100100111010000    0100100111010001    0100100111010010    0100100111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18895 - 18899

  --0100100111010100    0100100111010101    0100100111010110    0100100111010111    0100100111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18900 - 18904

  --0100100111011001    0100100111011010    0100100111011011    0100100111011100    0100100111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18905 - 18909

  --0100100111011110    0100100111011111    0100100111100000    0100100111100001    0100100111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18910 - 18914

  --0100100111100011    0100100111100100    0100100111100101    0100100111100110    0100100111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18915 - 18919

  --0100100111101000    0100100111101001    0100100111101010    0100100111101011    0100100111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18920 - 18924

  --0100100111101101    0100100111101110    0100100111101111    0100100111110000    0100100111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18925 - 18929

  --0100100111110010    0100100111110011    0100100111110100    0100100111110101    0100100111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18930 - 18934

  --0100100111110111    0100100111111000    0100100111111001    0100100111111010    0100100111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18935 - 18939

  --0100100111111100    0100100111111101    0100100111111110    0100100111111111    0100101000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18940 - 18944

  --0100101000000001    0100101000000010    0100101000000011    0100101000000100    0100101000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18945 - 18949

  --0100101000000110    0100101000000111    0100101000001000    0100101000001001    0100101000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18950 - 18954

  --0100101000001011    0100101000001100    0100101000001101    0100101000001110    0100101000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18955 - 18959

  --0100101000010000    0100101000010001    0100101000010010    0100101000010011    0100101000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18960 - 18964

  --0100101000010101    0100101000010110    0100101000010111    0100101000011000    0100101000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18965 - 18969

  --0100101000011010    0100101000011011    0100101000011100    0100101000011101    0100101000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18970 - 18974

  --0100101000011111    0100101000100000    0100101000100001    0100101000100010    0100101000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18975 - 18979

  --0100101000100100    0100101000100101    0100101000100110    0100101000100111    0100101000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18980 - 18984

  --0100101000101001    0100101000101010    0100101000101011    0100101000101100    0100101000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18985 - 18989

  --0100101000101110    0100101000101111    0100101000110000    0100101000110001    0100101000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18990 - 18994

  --0100101000110011    0100101000110100    0100101000110101    0100101000110110    0100101000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 18995 - 18999

  --0100101000111000    0100101000111001    0100101000111010    0100101000111011    0100101000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19000 - 19004

  --0100101000111101    0100101000111110    0100101000111111    0100101001000000    0100101001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19005 - 19009

  --0100101001000010    0100101001000011    0100101001000100    0100101001000101    0100101001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19010 - 19014

  --0100101001000111    0100101001001000    0100101001001001    0100101001001010    0100101001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19015 - 19019

  --0100101001001100    0100101001001101    0100101001001110    0100101001001111    0100101001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19020 - 19024

  --0100101001010001    0100101001010010    0100101001010011    0100101001010100    0100101001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19025 - 19029

  --0100101001010110    0100101001010111    0100101001011000    0100101001011001    0100101001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19030 - 19034

  --0100101001011011    0100101001011100    0100101001011101    0100101001011110    0100101001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19035 - 19039

  --0100101001100000    0100101001100001    0100101001100010    0100101001100011    0100101001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19040 - 19044

  --0100101001100101    0100101001100110    0100101001100111    0100101001101000    0100101001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19045 - 19049

  --0100101001101010    0100101001101011    0100101001101100    0100101001101101    0100101001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19050 - 19054

  --0100101001101111    0100101001110000    0100101001110001    0100101001110010    0100101001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19055 - 19059

  --0100101001110100    0100101001110101    0100101001110110    0100101001110111    0100101001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19060 - 19064

  --0100101001111001    0100101001111010    0100101001111011    0100101001111100    0100101001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19065 - 19069

  --0100101001111110    0100101001111111    0100101010000000    0100101010000001    0100101010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19070 - 19074

  --0100101010000011    0100101010000100    0100101010000101    0100101010000110    0100101010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19075 - 19079

  --0100101010001000    0100101010001001    0100101010001010    0100101010001011    0100101010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19080 - 19084

  --0100101010001101    0100101010001110    0100101010001111    0100101010010000    0100101010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19085 - 19089

  --0100101010010010    0100101010010011    0100101010010100    0100101010010101    0100101010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19090 - 19094

  --0100101010010111    0100101010011000    0100101010011001    0100101010011010    0100101010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19095 - 19099

  --0100101010011100    0100101010011101    0100101010011110    0100101010011111    0100101010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19100 - 19104

  --0100101010100001    0100101010100010    0100101010100011    0100101010100100    0100101010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19105 - 19109

  --0100101010100110    0100101010100111    0100101010101000    0100101010101001    0100101010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19110 - 19114

  --0100101010101011    0100101010101100    0100101010101101    0100101010101110    0100101010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19115 - 19119

  --0100101010110000    0100101010110001    0100101010110010    0100101010110011    0100101010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19120 - 19124

  --0100101010110101    0100101010110110    0100101010110111    0100101010111000    0100101010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19125 - 19129

  --0100101010111010    0100101010111011    0100101010111100    0100101010111101    0100101010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19130 - 19134

  --0100101010111111    0100101011000000    0100101011000001    0100101011000010    0100101011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19135 - 19139

  --0100101011000100    0100101011000101    0100101011000110    0100101011000111    0100101011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19140 - 19144

  --0100101011001001    0100101011001010    0100101011001011    0100101011001100    0100101011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19145 - 19149

  --0100101011001110    0100101011001111    0100101011010000    0100101011010001    0100101011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19150 - 19154

  --0100101011010011    0100101011010100    0100101011010101    0100101011010110    0100101011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19155 - 19159

  --0100101011011000    0100101011011001    0100101011011010    0100101011011011    0100101011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19160 - 19164

  --0100101011011101    0100101011011110    0100101011011111    0100101011100000    0100101011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19165 - 19169

  --0100101011100010    0100101011100011    0100101011100100    0100101011100101    0100101011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19170 - 19174

  --0100101011100111    0100101011101000    0100101011101001    0100101011101010    0100101011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19175 - 19179

  --0100101011101100    0100101011101101    0100101011101110    0100101011101111    0100101011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19180 - 19184

  --0100101011110001    0100101011110010    0100101011110011    0100101011110100    0100101011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19185 - 19189

  --0100101011110110    0100101011110111    0100101011111000    0100101011111001    0100101011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19190 - 19194

  --0100101011111011    0100101011111100    0100101011111101    0100101011111110    0100101011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19195 - 19199

  --0100101100000000    0100101100000001    0100101100000010    0100101100000011    0100101100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19200 - 19204

  --0100101100000101    0100101100000110    0100101100000111    0100101100001000    0100101100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19205 - 19209

  --0100101100001010    0100101100001011    0100101100001100    0100101100001101    0100101100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19210 - 19214

  --0100101100001111    0100101100010000    0100101100010001    0100101100010010    0100101100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19215 - 19219

  --0100101100010100    0100101100010101    0100101100010110    0100101100010111    0100101100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19220 - 19224

  --0100101100011001    0100101100011010    0100101100011011    0100101100011100    0100101100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19225 - 19229

  --0100101100011110    0100101100011111    0100101100100000    0100101100100001    0100101100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19230 - 19234

  --0100101100100011    0100101100100100    0100101100100101    0100101100100110    0100101100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19235 - 19239

  --0100101100101000    0100101100101001    0100101100101010    0100101100101011    0100101100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19240 - 19244

  --0100101100101101    0100101100101110    0100101100101111    0100101100110000    0100101100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19245 - 19249

  --0100101100110010    0100101100110011    0100101100110100    0100101100110101    0100101100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19250 - 19254

  --0100101100110111    0100101100111000    0100101100111001    0100101100111010    0100101100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19255 - 19259

  --0100101100111100    0100101100111101    0100101100111110    0100101100111111    0100101101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19260 - 19264

  --0100101101000001    0100101101000010    0100101101000011    0100101101000100    0100101101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19265 - 19269

  --0100101101000110    0100101101000111    0100101101001000    0100101101001001    0100101101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19270 - 19274

  --0100101101001011    0100101101001100    0100101101001101    0100101101001110    0100101101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19275 - 19279

  --0100101101010000    0100101101010001    0100101101010010    0100101101010011    0100101101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19280 - 19284

  --0100101101010101    0100101101010110    0100101101010111    0100101101011000    0100101101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19285 - 19289

  --0100101101011010    0100101101011011    0100101101011100    0100101101011101    0100101101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19290 - 19294

  --0100101101011111    0100101101100000    0100101101100001    0100101101100010    0100101101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19295 - 19299

  --0100101101100100    0100101101100101    0100101101100110    0100101101100111    0100101101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19300 - 19304

  --0100101101101001    0100101101101010    0100101101101011    0100101101101100    0100101101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19305 - 19309

  --0100101101101110    0100101101101111    0100101101110000    0100101101110001    0100101101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19310 - 19314

  --0100101101110011    0100101101110100    0100101101110101    0100101101110110    0100101101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19315 - 19319

  --0100101101111000    0100101101111001    0100101101111010    0100101101111011    0100101101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19320 - 19324

  --0100101101111101    0100101101111110    0100101101111111    0100101110000000    0100101110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19325 - 19329

  --0100101110000010    0100101110000011    0100101110000100    0100101110000101    0100101110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19330 - 19334

  --0100101110000111    0100101110001000    0100101110001001    0100101110001010    0100101110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19335 - 19339

  --0100101110001100    0100101110001101    0100101110001110    0100101110001111    0100101110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19340 - 19344

  --0100101110010001    0100101110010010    0100101110010011    0100101110010100    0100101110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19345 - 19349

  --0100101110010110    0100101110010111    0100101110011000    0100101110011001    0100101110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19350 - 19354

  --0100101110011011    0100101110011100    0100101110011101    0100101110011110    0100101110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19355 - 19359

  --0100101110100000    0100101110100001    0100101110100010    0100101110100011    0100101110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19360 - 19364

  --0100101110100101    0100101110100110    0100101110100111    0100101110101000    0100101110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19365 - 19369

  --0100101110101010    0100101110101011    0100101110101100    0100101110101101    0100101110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19370 - 19374

  --0100101110101111    0100101110110000    0100101110110001    0100101110110010    0100101110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19375 - 19379

  --0100101110110100    0100101110110101    0100101110110110    0100101110110111    0100101110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19380 - 19384

  --0100101110111001    0100101110111010    0100101110111011    0100101110111100    0100101110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19385 - 19389

  --0100101110111110    0100101110111111    0100101111000000    0100101111000001    0100101111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19390 - 19394

  --0100101111000011    0100101111000100    0100101111000101    0100101111000110    0100101111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19395 - 19399

  --0100101111001000    0100101111001001    0100101111001010    0100101111001011    0100101111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19400 - 19404

  --0100101111001101    0100101111001110    0100101111001111    0100101111010000    0100101111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19405 - 19409

  --0100101111010010    0100101111010011    0100101111010100    0100101111010101    0100101111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19410 - 19414

  --0100101111010111    0100101111011000    0100101111011001    0100101111011010    0100101111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19415 - 19419

  --0100101111011100    0100101111011101    0100101111011110    0100101111011111    0100101111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19420 - 19424

  --0100101111100001    0100101111100010    0100101111100011    0100101111100100    0100101111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19425 - 19429

  --0100101111100110    0100101111100111    0100101111101000    0100101111101001    0100101111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19430 - 19434

  --0100101111101011    0100101111101100    0100101111101101    0100101111101110    0100101111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19435 - 19439

  --0100101111110000    0100101111110001    0100101111110010    0100101111110011    0100101111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19440 - 19444

  --0100101111110101    0100101111110110    0100101111110111    0100101111111000    0100101111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19445 - 19449

  --0100101111111010    0100101111111011    0100101111111100    0100101111111101    0100101111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19450 - 19454

  --0100101111111111    0100110000000000    0100110000000001    0100110000000010    0100110000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19455 - 19459

  --0100110000000100    0100110000000101    0100110000000110    0100110000000111    0100110000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19460 - 19464

  --0100110000001001    0100110000001010    0100110000001011    0100110000001100    0100110000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19465 - 19469

  --0100110000001110    0100110000001111    0100110000010000    0100110000010001    0100110000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19470 - 19474

  --0100110000010011    0100110000010100    0100110000010101    0100110000010110    0100110000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19475 - 19479

  --0100110000011000    0100110000011001    0100110000011010    0100110000011011    0100110000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19480 - 19484

  --0100110000011101    0100110000011110    0100110000011111    0100110000100000    0100110000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19485 - 19489

  --0100110000100010    0100110000100011    0100110000100100    0100110000100101    0100110000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19490 - 19494

  --0100110000100111    0100110000101000    0100110000101001    0100110000101010    0100110000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19495 - 19499

  --0100110000101100    0100110000101101    0100110000101110    0100110000101111    0100110000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19500 - 19504

  --0100110000110001    0100110000110010    0100110000110011    0100110000110100    0100110000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19505 - 19509

  --0100110000110110    0100110000110111    0100110000111000    0100110000111001    0100110000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19510 - 19514

  --0100110000111011    0100110000111100    0100110000111101    0100110000111110    0100110000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19515 - 19519

  --0100110001000000    0100110001000001    0100110001000010    0100110001000011    0100110001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19520 - 19524

  --0100110001000101    0100110001000110    0100110001000111    0100110001001000    0100110001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19525 - 19529

  --0100110001001010    0100110001001011    0100110001001100    0100110001001101    0100110001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19530 - 19534

  --0100110001001111    0100110001010000    0100110001010001    0100110001010010    0100110001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19535 - 19539

  --0100110001010100    0100110001010101    0100110001010110    0100110001010111    0100110001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19540 - 19544

  --0100110001011001    0100110001011010    0100110001011011    0100110001011100    0100110001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19545 - 19549

  --0100110001011110    0100110001011111    0100110001100000    0100110001100001    0100110001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19550 - 19554

  --0100110001100011    0100110001100100    0100110001100101    0100110001100110    0100110001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19555 - 19559

  --0100110001101000    0100110001101001    0100110001101010    0100110001101011    0100110001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19560 - 19564

  --0100110001101101    0100110001101110    0100110001101111    0100110001110000    0100110001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19565 - 19569

  --0100110001110010    0100110001110011    0100110001110100    0100110001110101    0100110001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19570 - 19574

  --0100110001110111    0100110001111000    0100110001111001    0100110001111010    0100110001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19575 - 19579

  --0100110001111100    0100110001111101    0100110001111110    0100110001111111    0100110010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19580 - 19584

  --0100110010000001    0100110010000010    0100110010000011    0100110010000100    0100110010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19585 - 19589

  --0100110010000110    0100110010000111    0100110010001000    0100110010001001    0100110010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19590 - 19594

  --0100110010001011    0100110010001100    0100110010001101    0100110010001110    0100110010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19595 - 19599

  --0100110010010000    0100110010010001    0100110010010010    0100110010010011    0100110010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19600 - 19604

  --0100110010010101    0100110010010110    0100110010010111    0100110010011000    0100110010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19605 - 19609

  --0100110010011010    0100110010011011    0100110010011100    0100110010011101    0100110010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19610 - 19614

  --0100110010011111    0100110010100000    0100110010100001    0100110010100010    0100110010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19615 - 19619

  --0100110010100100    0100110010100101    0100110010100110    0100110010100111    0100110010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19620 - 19624

  --0100110010101001    0100110010101010    0100110010101011    0100110010101100    0100110010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19625 - 19629

  --0100110010101110    0100110010101111    0100110010110000    0100110010110001    0100110010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19630 - 19634

  --0100110010110011    0100110010110100    0100110010110101    0100110010110110    0100110010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19635 - 19639

  --0100110010111000    0100110010111001    0100110010111010    0100110010111011    0100110010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19640 - 19644

  --0100110010111101    0100110010111110    0100110010111111    0100110011000000    0100110011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19645 - 19649

  --0100110011000010    0100110011000011    0100110011000100    0100110011000101    0100110011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19650 - 19654

  --0100110011000111    0100110011001000    0100110011001001    0100110011001010    0100110011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19655 - 19659

  --0100110011001100    0100110011001101    0100110011001110    0100110011001111    0100110011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19660 - 19664

  --0100110011010001    0100110011010010    0100110011010011    0100110011010100    0100110011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19665 - 19669

  --0100110011010110    0100110011010111    0100110011011000    0100110011011001    0100110011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19670 - 19674

  --0100110011011011    0100110011011100    0100110011011101    0100110011011110    0100110011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19675 - 19679

  --0100110011100000    0100110011100001    0100110011100010    0100110011100011    0100110011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19680 - 19684

  --0100110011100101    0100110011100110    0100110011100111    0100110011101000    0100110011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19685 - 19689

  --0100110011101010    0100110011101011    0100110011101100    0100110011101101    0100110011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19690 - 19694

  --0100110011101111    0100110011110000    0100110011110001    0100110011110010    0100110011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19695 - 19699

  --0100110011110100    0100110011110101    0100110011110110    0100110011110111    0100110011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19700 - 19704

  --0100110011111001    0100110011111010    0100110011111011    0100110011111100    0100110011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19705 - 19709

  --0100110011111110    0100110011111111    0100110100000000    0100110100000001    0100110100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19710 - 19714

  --0100110100000011    0100110100000100    0100110100000101    0100110100000110    0100110100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19715 - 19719

  --0100110100001000    0100110100001001    0100110100001010    0100110100001011    0100110100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19720 - 19724

  --0100110100001101    0100110100001110    0100110100001111    0100110100010000    0100110100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19725 - 19729

  --0100110100010010    0100110100010011    0100110100010100    0100110100010101    0100110100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19730 - 19734

  --0100110100010111    0100110100011000    0100110100011001    0100110100011010    0100110100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19735 - 19739

  --0100110100011100    0100110100011101    0100110100011110    0100110100011111    0100110100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19740 - 19744

  --0100110100100001    0100110100100010    0100110100100011    0100110100100100    0100110100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19745 - 19749

  --0100110100100110    0100110100100111    0100110100101000    0100110100101001    0100110100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19750 - 19754

  --0100110100101011    0100110100101100    0100110100101101    0100110100101110    0100110100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19755 - 19759

  --0100110100110000    0100110100110001    0100110100110010    0100110100110011    0100110100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19760 - 19764

  --0100110100110101    0100110100110110    0100110100110111    0100110100111000    0100110100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19765 - 19769

  --0100110100111010    0100110100111011    0100110100111100    0100110100111101    0100110100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19770 - 19774

  --0100110100111111    0100110101000000    0100110101000001    0100110101000010    0100110101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19775 - 19779

  --0100110101000100    0100110101000101    0100110101000110    0100110101000111    0100110101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19780 - 19784

  --0100110101001001    0100110101001010    0100110101001011    0100110101001100    0100110101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19785 - 19789

  --0100110101001110    0100110101001111    0100110101010000    0100110101010001    0100110101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19790 - 19794

  --0100110101010011    0100110101010100    0100110101010101    0100110101010110    0100110101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19795 - 19799

  --0100110101011000    0100110101011001    0100110101011010    0100110101011011    0100110101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19800 - 19804

  --0100110101011101    0100110101011110    0100110101011111    0100110101100000    0100110101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19805 - 19809

  --0100110101100010    0100110101100011    0100110101100100    0100110101100101    0100110101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19810 - 19814

  --0100110101100111    0100110101101000    0100110101101001    0100110101101010    0100110101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19815 - 19819

  --0100110101101100    0100110101101101    0100110101101110    0100110101101111    0100110101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19820 - 19824

  --0100110101110001    0100110101110010    0100110101110011    0100110101110100    0100110101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19825 - 19829

  --0100110101110110    0100110101110111    0100110101111000    0100110101111001    0100110101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19830 - 19834

  --0100110101111011    0100110101111100    0100110101111101    0100110101111110    0100110101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19835 - 19839

  --0100110110000000    0100110110000001    0100110110000010    0100110110000011    0100110110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19840 - 19844

  --0100110110000101    0100110110000110    0100110110000111    0100110110001000    0100110110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19845 - 19849

  --0100110110001010    0100110110001011    0100110110001100    0100110110001101    0100110110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19850 - 19854

  --0100110110001111    0100110110010000    0100110110010001    0100110110010010    0100110110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19855 - 19859

  --0100110110010100    0100110110010101    0100110110010110    0100110110010111    0100110110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19860 - 19864

  --0100110110011001    0100110110011010    0100110110011011    0100110110011100    0100110110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19865 - 19869

  --0100110110011110    0100110110011111    0100110110100000    0100110110100001    0100110110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19870 - 19874

  --0100110110100011    0100110110100100    0100110110100101    0100110110100110    0100110110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19875 - 19879

  --0100110110101000    0100110110101001    0100110110101010    0100110110101011    0100110110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19880 - 19884

  --0100110110101101    0100110110101110    0100110110101111    0100110110110000    0100110110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19885 - 19889

  --0100110110110010    0100110110110011    0100110110110100    0100110110110101    0100110110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19890 - 19894

  --0100110110110111    0100110110111000    0100110110111001    0100110110111010    0100110110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19895 - 19899

  --0100110110111100    0100110110111101    0100110110111110    0100110110111111    0100110111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19900 - 19904

  --0100110111000001    0100110111000010    0100110111000011    0100110111000100    0100110111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19905 - 19909

  --0100110111000110    0100110111000111    0100110111001000    0100110111001001    0100110111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19910 - 19914

  --0100110111001011    0100110111001100    0100110111001101    0100110111001110    0100110111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19915 - 19919

  --0100110111010000    0100110111010001    0100110111010010    0100110111010011    0100110111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19920 - 19924

  --0100110111010101    0100110111010110    0100110111010111    0100110111011000    0100110111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19925 - 19929

  --0100110111011010    0100110111011011    0100110111011100    0100110111011101    0100110111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19930 - 19934

  --0100110111011111    0100110111100000    0100110111100001    0100110111100010    0100110111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19935 - 19939

  --0100110111100100    0100110111100101    0100110111100110    0100110111100111    0100110111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19940 - 19944

  --0100110111101001    0100110111101010    0100110111101011    0100110111101100    0100110111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19945 - 19949

  --0100110111101110    0100110111101111    0100110111110000    0100110111110001    0100110111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19950 - 19954

  --0100110111110011    0100110111110100    0100110111110101    0100110111110110    0100110111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19955 - 19959

  --0100110111111000    0100110111111001    0100110111111010    0100110111111011    0100110111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19960 - 19964

  --0100110111111101    0100110111111110    0100110111111111    0100111000000000    0100111000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19965 - 19969

  --0100111000000010    0100111000000011    0100111000000100    0100111000000101    0100111000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19970 - 19974

  --0100111000000111    0100111000001000    0100111000001001    0100111000001010    0100111000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19975 - 19979

  --0100111000001100    0100111000001101    0100111000001110    0100111000001111    0100111000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19980 - 19984

  --0100111000010001    0100111000010010    0100111000010011    0100111000010100    0100111000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19985 - 19989

  --0100111000010110    0100111000010111    0100111000011000    0100111000011001    0100111000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19990 - 19994

  --0100111000011011    0100111000011100    0100111000011101    0100111000011110    0100111000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 19995 - 19999

  --0100111000100000    0100111000100001    0100111000100010    0100111000100011    0100111000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20000 - 20004

  --0100111000100101    0100111000100110    0100111000100111    0100111000101000    0100111000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20005 - 20009

  --0100111000101010    0100111000101011    0100111000101100    0100111000101101    0100111000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20010 - 20014

  --0100111000101111    0100111000110000    0100111000110001    0100111000110010    0100111000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20015 - 20019

  --0100111000110100    0100111000110101    0100111000110110    0100111000110111    0100111000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20020 - 20024

  --0100111000111001    0100111000111010    0100111000111011    0100111000111100    0100111000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20025 - 20029

  --0100111000111110    0100111000111111    0100111001000000    0100111001000001    0100111001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20030 - 20034

  --0100111001000011    0100111001000100    0100111001000101    0100111001000110    0100111001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20035 - 20039

  --0100111001001000    0100111001001001    0100111001001010    0100111001001011    0100111001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20040 - 20044

  --0100111001001101    0100111001001110    0100111001001111    0100111001010000    0100111001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20045 - 20049

  --0100111001010010    0100111001010011    0100111001010100    0100111001010101    0100111001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20050 - 20054

  --0100111001010111    0100111001011000    0100111001011001    0100111001011010    0100111001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20055 - 20059

  --0100111001011100    0100111001011101    0100111001011110    0100111001011111    0100111001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20060 - 20064

  --0100111001100001    0100111001100010    0100111001100011    0100111001100100    0100111001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20065 - 20069

  --0100111001100110    0100111001100111    0100111001101000    0100111001101001    0100111001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20070 - 20074

  --0100111001101011    0100111001101100    0100111001101101    0100111001101110    0100111001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20075 - 20079

  --0100111001110000    0100111001110001    0100111001110010    0100111001110011    0100111001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20080 - 20084

  --0100111001110101    0100111001110110    0100111001110111    0100111001111000    0100111001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20085 - 20089

  --0100111001111010    0100111001111011    0100111001111100    0100111001111101    0100111001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20090 - 20094

  --0100111001111111    0100111010000000    0100111010000001    0100111010000010    0100111010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20095 - 20099

  --0100111010000100    0100111010000101    0100111010000110    0100111010000111    0100111010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20100 - 20104

  --0100111010001001    0100111010001010    0100111010001011    0100111010001100    0100111010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20105 - 20109

  --0100111010001110    0100111010001111    0100111010010000    0100111010010001    0100111010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20110 - 20114

  --0100111010010011    0100111010010100    0100111010010101    0100111010010110    0100111010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20115 - 20119

  --0100111010011000    0100111010011001    0100111010011010    0100111010011011    0100111010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20120 - 20124

  --0100111010011101    0100111010011110    0100111010011111    0100111010100000    0100111010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20125 - 20129

  --0100111010100010    0100111010100011    0100111010100100    0100111010100101    0100111010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20130 - 20134

  --0100111010100111    0100111010101000    0100111010101001    0100111010101010    0100111010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20135 - 20139

  --0100111010101100    0100111010101101    0100111010101110    0100111010101111    0100111010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20140 - 20144

  --0100111010110001    0100111010110010    0100111010110011    0100111010110100    0100111010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20145 - 20149

  --0100111010110110    0100111010110111    0100111010111000    0100111010111001    0100111010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20150 - 20154

  --0100111010111011    0100111010111100    0100111010111101    0100111010111110    0100111010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20155 - 20159

  --0100111011000000    0100111011000001    0100111011000010    0100111011000011    0100111011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20160 - 20164

  --0100111011000101    0100111011000110    0100111011000111    0100111011001000    0100111011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20165 - 20169

  --0100111011001010    0100111011001011    0100111011001100    0100111011001101    0100111011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20170 - 20174

  --0100111011001111    0100111011010000    0100111011010001    0100111011010010    0100111011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20175 - 20179

  --0100111011010100    0100111011010101    0100111011010110    0100111011010111    0100111011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20180 - 20184

  --0100111011011001    0100111011011010    0100111011011011    0100111011011100    0100111011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20185 - 20189

  --0100111011011110    0100111011011111    0100111011100000    0100111011100001    0100111011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20190 - 20194

  --0100111011100011    0100111011100100    0100111011100101    0100111011100110    0100111011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20195 - 20199

  --0100111011101000    0100111011101001    0100111011101010    0100111011101011    0100111011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20200 - 20204

  --0100111011101101    0100111011101110    0100111011101111    0100111011110000    0100111011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20205 - 20209

  --0100111011110010    0100111011110011    0100111011110100    0100111011110101    0100111011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20210 - 20214

  --0100111011110111    0100111011111000    0100111011111001    0100111011111010    0100111011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20215 - 20219

  --0100111011111100    0100111011111101    0100111011111110    0100111011111111    0100111100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20220 - 20224

  --0100111100000001    0100111100000010    0100111100000011    0100111100000100    0100111100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20225 - 20229

  --0100111100000110    0100111100000111    0100111100001000    0100111100001001    0100111100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20230 - 20234

  --0100111100001011    0100111100001100    0100111100001101    0100111100001110    0100111100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20235 - 20239

  --0100111100010000    0100111100010001    0100111100010010    0100111100010011    0100111100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20240 - 20244

  --0100111100010101    0100111100010110    0100111100010111    0100111100011000    0100111100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20245 - 20249

  --0100111100011010    0100111100011011    0100111100011100    0100111100011101    0100111100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20250 - 20254

  --0100111100011111    0100111100100000    0100111100100001    0100111100100010    0100111100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20255 - 20259

  --0100111100100100    0100111100100101    0100111100100110    0100111100100111    0100111100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20260 - 20264

  --0100111100101001    0100111100101010    0100111100101011    0100111100101100    0100111100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20265 - 20269

  --0100111100101110    0100111100101111    0100111100110000    0100111100110001    0100111100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20270 - 20274

  --0100111100110011    0100111100110100    0100111100110101    0100111100110110    0100111100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20275 - 20279

  --0100111100111000    0100111100111001    0100111100111010    0100111100111011    0100111100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20280 - 20284

  --0100111100111101    0100111100111110    0100111100111111    0100111101000000    0100111101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20285 - 20289

  --0100111101000010    0100111101000011    0100111101000100    0100111101000101    0100111101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20290 - 20294

  --0100111101000111    0100111101001000    0100111101001001    0100111101001010    0100111101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20295 - 20299

  --0100111101001100    0100111101001101    0100111101001110    0100111101001111    0100111101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20300 - 20304

  --0100111101010001    0100111101010010    0100111101010011    0100111101010100    0100111101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20305 - 20309

  --0100111101010110    0100111101010111    0100111101011000    0100111101011001    0100111101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20310 - 20314

  --0100111101011011    0100111101011100    0100111101011101    0100111101011110    0100111101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20315 - 20319

  --0100111101100000    0100111101100001    0100111101100010    0100111101100011    0100111101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20320 - 20324

  --0100111101100101    0100111101100110    0100111101100111    0100111101101000    0100111101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20325 - 20329

  --0100111101101010    0100111101101011    0100111101101100    0100111101101101    0100111101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20330 - 20334

  --0100111101101111    0100111101110000    0100111101110001    0100111101110010    0100111101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20335 - 20339

  --0100111101110100    0100111101110101    0100111101110110    0100111101110111    0100111101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20340 - 20344

  --0100111101111001    0100111101111010    0100111101111011    0100111101111100    0100111101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20345 - 20349

  --0100111101111110    0100111101111111    0100111110000000    0100111110000001    0100111110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20350 - 20354

  --0100111110000011    0100111110000100    0100111110000101    0100111110000110    0100111110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20355 - 20359

  --0100111110001000    0100111110001001    0100111110001010    0100111110001011    0100111110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20360 - 20364

  --0100111110001101    0100111110001110    0100111110001111    0100111110010000    0100111110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20365 - 20369

  --0100111110010010    0100111110010011    0100111110010100    0100111110010101    0100111110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20370 - 20374

  --0100111110010111    0100111110011000    0100111110011001    0100111110011010    0100111110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20375 - 20379

  --0100111110011100    0100111110011101    0100111110011110    0100111110011111    0100111110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20380 - 20384

  --0100111110100001    0100111110100010    0100111110100011    0100111110100100    0100111110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20385 - 20389

  --0100111110100110    0100111110100111    0100111110101000    0100111110101001    0100111110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20390 - 20394

  --0100111110101011    0100111110101100    0100111110101101    0100111110101110    0100111110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20395 - 20399

  --0100111110110000    0100111110110001    0100111110110010    0100111110110011    0100111110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20400 - 20404

  --0100111110110101    0100111110110110    0100111110110111    0100111110111000    0100111110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20405 - 20409

  --0100111110111010    0100111110111011    0100111110111100    0100111110111101    0100111110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20410 - 20414

  --0100111110111111    0100111111000000    0100111111000001    0100111111000010    0100111111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20415 - 20419

  --0100111111000100    0100111111000101    0100111111000110    0100111111000111    0100111111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20420 - 20424

  --0100111111001001    0100111111001010    0100111111001011    0100111111001100    0100111111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20425 - 20429

  --0100111111001110    0100111111001111    0100111111010000    0100111111010001    0100111111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20430 - 20434

  --0100111111010011    0100111111010100    0100111111010101    0100111111010110    0100111111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20435 - 20439

  --0100111111011000    0100111111011001    0100111111011010    0100111111011011    0100111111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20440 - 20444

  --0100111111011101    0100111111011110    0100111111011111    0100111111100000    0100111111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20445 - 20449

  --0100111111100010    0100111111100011    0100111111100100    0100111111100101    0100111111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20450 - 20454

  --0100111111100111    0100111111101000    0100111111101001    0100111111101010    0100111111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20455 - 20459

  --0100111111101100    0100111111101101    0100111111101110    0100111111101111    0100111111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20460 - 20464

  --0100111111110001    0100111111110010    0100111111110011    0100111111110100    0100111111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20465 - 20469

  --0100111111110110    0100111111110111    0100111111111000    0100111111111001    0100111111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20470 - 20474

  --0100111111111011    0100111111111100    0100111111111101    0100111111111110    0100111111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20475 - 20479

  --0101000000000000    0101000000000001    0101000000000010    0101000000000011    0101000000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20480 - 20484

  --0101000000000101    0101000000000110    0101000000000111    0101000000001000    0101000000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20485 - 20489

  --0101000000001010    0101000000001011    0101000000001100    0101000000001101    0101000000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20490 - 20494

  --0101000000001111    0101000000010000    0101000000010001    0101000000010010    0101000000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20495 - 20499

  --0101000000010100    0101000000010101    0101000000010110    0101000000010111    0101000000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20500 - 20504

  --0101000000011001    0101000000011010    0101000000011011    0101000000011100    0101000000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20505 - 20509

  --0101000000011110    0101000000011111    0101000000100000    0101000000100001    0101000000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20510 - 20514

  --0101000000100011    0101000000100100    0101000000100101    0101000000100110    0101000000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20515 - 20519

  --0101000000101000    0101000000101001    0101000000101010    0101000000101011    0101000000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20520 - 20524

  --0101000000101101    0101000000101110    0101000000101111    0101000000110000    0101000000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20525 - 20529

  --0101000000110010    0101000000110011    0101000000110100    0101000000110101    0101000000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20530 - 20534

  --0101000000110111    0101000000111000    0101000000111001    0101000000111010    0101000000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20535 - 20539

  --0101000000111100    0101000000111101    0101000000111110    0101000000111111    0101000001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20540 - 20544

  --0101000001000001    0101000001000010    0101000001000011    0101000001000100    0101000001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20545 - 20549

  --0101000001000110    0101000001000111    0101000001001000    0101000001001001    0101000001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20550 - 20554

  --0101000001001011    0101000001001100    0101000001001101    0101000001001110    0101000001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20555 - 20559

  --0101000001010000    0101000001010001    0101000001010010    0101000001010011    0101000001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20560 - 20564

  --0101000001010101    0101000001010110    0101000001010111    0101000001011000    0101000001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20565 - 20569

  --0101000001011010    0101000001011011    0101000001011100    0101000001011101    0101000001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20570 - 20574

  --0101000001011111    0101000001100000    0101000001100001    0101000001100010    0101000001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20575 - 20579

  --0101000001100100    0101000001100101    0101000001100110    0101000001100111    0101000001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20580 - 20584

  --0101000001101001    0101000001101010    0101000001101011    0101000001101100    0101000001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20585 - 20589

  --0101000001101110    0101000001101111    0101000001110000    0101000001110001    0101000001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20590 - 20594

  --0101000001110011    0101000001110100    0101000001110101    0101000001110110    0101000001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20595 - 20599

  --0101000001111000    0101000001111001    0101000001111010    0101000001111011    0101000001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20600 - 20604

  --0101000001111101    0101000001111110    0101000001111111    0101000010000000    0101000010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20605 - 20609

  --0101000010000010    0101000010000011    0101000010000100    0101000010000101    0101000010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20610 - 20614

  --0101000010000111    0101000010001000    0101000010001001    0101000010001010    0101000010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20615 - 20619

  --0101000010001100    0101000010001101    0101000010001110    0101000010001111    0101000010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20620 - 20624

  --0101000010010001    0101000010010010    0101000010010011    0101000010010100    0101000010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20625 - 20629

  --0101000010010110    0101000010010111    0101000010011000    0101000010011001    0101000010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20630 - 20634

  --0101000010011011    0101000010011100    0101000010011101    0101000010011110    0101000010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20635 - 20639

  --0101000010100000    0101000010100001    0101000010100010    0101000010100011    0101000010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20640 - 20644

  --0101000010100101    0101000010100110    0101000010100111    0101000010101000    0101000010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20645 - 20649

  --0101000010101010    0101000010101011    0101000010101100    0101000010101101    0101000010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20650 - 20654

  --0101000010101111    0101000010110000    0101000010110001    0101000010110010    0101000010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20655 - 20659

  --0101000010110100    0101000010110101    0101000010110110    0101000010110111    0101000010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20660 - 20664

  --0101000010111001    0101000010111010    0101000010111011    0101000010111100    0101000010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20665 - 20669

  --0101000010111110    0101000010111111    0101000011000000    0101000011000001    0101000011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20670 - 20674

  --0101000011000011    0101000011000100    0101000011000101    0101000011000110    0101000011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20675 - 20679

  --0101000011001000    0101000011001001    0101000011001010    0101000011001011    0101000011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20680 - 20684

  --0101000011001101    0101000011001110    0101000011001111    0101000011010000    0101000011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20685 - 20689

  --0101000011010010    0101000011010011    0101000011010100    0101000011010101    0101000011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20690 - 20694

  --0101000011010111    0101000011011000    0101000011011001    0101000011011010    0101000011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20695 - 20699

  --0101000011011100    0101000011011101    0101000011011110    0101000011011111    0101000011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20700 - 20704

  --0101000011100001    0101000011100010    0101000011100011    0101000011100100    0101000011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20705 - 20709

  --0101000011100110    0101000011100111    0101000011101000    0101000011101001    0101000011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20710 - 20714

  --0101000011101011    0101000011101100    0101000011101101    0101000011101110    0101000011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20715 - 20719

  --0101000011110000    0101000011110001    0101000011110010    0101000011110011    0101000011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20720 - 20724

  --0101000011110101    0101000011110110    0101000011110111    0101000011111000    0101000011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20725 - 20729

  --0101000011111010    0101000011111011    0101000011111100    0101000011111101    0101000011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20730 - 20734

  --0101000011111111    0101000100000000    0101000100000001    0101000100000010    0101000100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20735 - 20739

  --0101000100000100    0101000100000101    0101000100000110    0101000100000111    0101000100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20740 - 20744

  --0101000100001001    0101000100001010    0101000100001011    0101000100001100    0101000100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20745 - 20749

  --0101000100001110    0101000100001111    0101000100010000    0101000100010001    0101000100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20750 - 20754

  --0101000100010011    0101000100010100    0101000100010101    0101000100010110    0101000100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20755 - 20759

  --0101000100011000    0101000100011001    0101000100011010    0101000100011011    0101000100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20760 - 20764

  --0101000100011101    0101000100011110    0101000100011111    0101000100100000    0101000100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20765 - 20769

  --0101000100100010    0101000100100011    0101000100100100    0101000100100101    0101000100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20770 - 20774

  --0101000100100111    0101000100101000    0101000100101001    0101000100101010    0101000100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20775 - 20779

  --0101000100101100    0101000100101101    0101000100101110    0101000100101111    0101000100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20780 - 20784

  --0101000100110001    0101000100110010    0101000100110011    0101000100110100    0101000100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20785 - 20789

  --0101000100110110    0101000100110111    0101000100111000    0101000100111001    0101000100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20790 - 20794

  --0101000100111011    0101000100111100    0101000100111101    0101000100111110    0101000100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20795 - 20799

  --0101000101000000    0101000101000001    0101000101000010    0101000101000011    0101000101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20800 - 20804

  --0101000101000101    0101000101000110    0101000101000111    0101000101001000    0101000101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20805 - 20809

  --0101000101001010    0101000101001011    0101000101001100    0101000101001101    0101000101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20810 - 20814

  --0101000101001111    0101000101010000    0101000101010001    0101000101010010    0101000101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20815 - 20819

  --0101000101010100    0101000101010101    0101000101010110    0101000101010111    0101000101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20820 - 20824

  --0101000101011001    0101000101011010    0101000101011011    0101000101011100    0101000101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20825 - 20829

  --0101000101011110    0101000101011111    0101000101100000    0101000101100001    0101000101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20830 - 20834

  --0101000101100011    0101000101100100    0101000101100101    0101000101100110    0101000101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20835 - 20839

  --0101000101101000    0101000101101001    0101000101101010    0101000101101011    0101000101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20840 - 20844

  --0101000101101101    0101000101101110    0101000101101111    0101000101110000    0101000101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20845 - 20849

  --0101000101110010    0101000101110011    0101000101110100    0101000101110101    0101000101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20850 - 20854

  --0101000101110111    0101000101111000    0101000101111001    0101000101111010    0101000101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20855 - 20859

  --0101000101111100    0101000101111101    0101000101111110    0101000101111111    0101000110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20860 - 20864

  --0101000110000001    0101000110000010    0101000110000011    0101000110000100    0101000110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20865 - 20869

  --0101000110000110    0101000110000111    0101000110001000    0101000110001001    0101000110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20870 - 20874

  --0101000110001011    0101000110001100    0101000110001101    0101000110001110    0101000110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20875 - 20879

  --0101000110010000    0101000110010001    0101000110010010    0101000110010011    0101000110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20880 - 20884

  --0101000110010101    0101000110010110    0101000110010111    0101000110011000    0101000110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20885 - 20889

  --0101000110011010    0101000110011011    0101000110011100    0101000110011101    0101000110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20890 - 20894

  --0101000110011111    0101000110100000    0101000110100001    0101000110100010    0101000110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20895 - 20899

  --0101000110100100    0101000110100101    0101000110100110    0101000110100111    0101000110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20900 - 20904

  --0101000110101001    0101000110101010    0101000110101011    0101000110101100    0101000110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20905 - 20909

  --0101000110101110    0101000110101111    0101000110110000    0101000110110001    0101000110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20910 - 20914

  --0101000110110011    0101000110110100    0101000110110101    0101000110110110    0101000110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20915 - 20919

  --0101000110111000    0101000110111001    0101000110111010    0101000110111011    0101000110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20920 - 20924

  --0101000110111101    0101000110111110    0101000110111111    0101000111000000    0101000111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20925 - 20929

  --0101000111000010    0101000111000011    0101000111000100    0101000111000101    0101000111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20930 - 20934

  --0101000111000111    0101000111001000    0101000111001001    0101000111001010    0101000111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20935 - 20939

  --0101000111001100    0101000111001101    0101000111001110    0101000111001111    0101000111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20940 - 20944

  --0101000111010001    0101000111010010    0101000111010011    0101000111010100    0101000111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20945 - 20949

  --0101000111010110    0101000111010111    0101000111011000    0101000111011001    0101000111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20950 - 20954

  --0101000111011011    0101000111011100    0101000111011101    0101000111011110    0101000111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20955 - 20959

  --0101000111100000    0101000111100001    0101000111100010    0101000111100011    0101000111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20960 - 20964

  --0101000111100101    0101000111100110    0101000111100111    0101000111101000    0101000111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20965 - 20969

  --0101000111101010    0101000111101011    0101000111101100    0101000111101101    0101000111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20970 - 20974

  --0101000111101111    0101000111110000    0101000111110001    0101000111110010    0101000111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20975 - 20979

  --0101000111110100    0101000111110101    0101000111110110    0101000111110111    0101000111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20980 - 20984

  --0101000111111001    0101000111111010    0101000111111011    0101000111111100    0101000111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20985 - 20989

  --0101000111111110    0101000111111111    0101001000000000    0101001000000001    0101001000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20990 - 20994

  --0101001000000011    0101001000000100    0101001000000101    0101001000000110    0101001000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 20995 - 20999

  --0101001000001000    0101001000001001    0101001000001010    0101001000001011    0101001000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21000 - 21004

  --0101001000001101    0101001000001110    0101001000001111    0101001000010000    0101001000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21005 - 21009

  --0101001000010010    0101001000010011    0101001000010100    0101001000010101    0101001000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21010 - 21014

  --0101001000010111    0101001000011000    0101001000011001    0101001000011010    0101001000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21015 - 21019

  --0101001000011100    0101001000011101    0101001000011110    0101001000011111    0101001000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21020 - 21024

  --0101001000100001    0101001000100010    0101001000100011    0101001000100100    0101001000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21025 - 21029

  --0101001000100110    0101001000100111    0101001000101000    0101001000101001    0101001000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21030 - 21034

  --0101001000101011    0101001000101100    0101001000101101    0101001000101110    0101001000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21035 - 21039

  --0101001000110000    0101001000110001    0101001000110010    0101001000110011    0101001000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21040 - 21044

  --0101001000110101    0101001000110110    0101001000110111    0101001000111000    0101001000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21045 - 21049

  --0101001000111010    0101001000111011    0101001000111100    0101001000111101    0101001000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21050 - 21054

  --0101001000111111    0101001001000000    0101001001000001    0101001001000010    0101001001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21055 - 21059

  --0101001001000100    0101001001000101    0101001001000110    0101001001000111    0101001001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21060 - 21064

  --0101001001001001    0101001001001010    0101001001001011    0101001001001100    0101001001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21065 - 21069

  --0101001001001110    0101001001001111    0101001001010000    0101001001010001    0101001001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21070 - 21074

  --0101001001010011    0101001001010100    0101001001010101    0101001001010110    0101001001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21075 - 21079

  --0101001001011000    0101001001011001    0101001001011010    0101001001011011    0101001001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21080 - 21084

  --0101001001011101    0101001001011110    0101001001011111    0101001001100000    0101001001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21085 - 21089

  --0101001001100010    0101001001100011    0101001001100100    0101001001100101    0101001001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21090 - 21094

  --0101001001100111    0101001001101000    0101001001101001    0101001001101010    0101001001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21095 - 21099

  --0101001001101100    0101001001101101    0101001001101110    0101001001101111    0101001001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21100 - 21104

  --0101001001110001    0101001001110010    0101001001110011    0101001001110100    0101001001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21105 - 21109

  --0101001001110110    0101001001110111    0101001001111000    0101001001111001    0101001001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21110 - 21114

  --0101001001111011    0101001001111100    0101001001111101    0101001001111110    0101001001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21115 - 21119

  --0101001010000000    0101001010000001    0101001010000010    0101001010000011    0101001010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21120 - 21124

  --0101001010000101    0101001010000110    0101001010000111    0101001010001000    0101001010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21125 - 21129

  --0101001010001010    0101001010001011    0101001010001100    0101001010001101    0101001010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21130 - 21134

  --0101001010001111    0101001010010000    0101001010010001    0101001010010010    0101001010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21135 - 21139

  --0101001010010100    0101001010010101    0101001010010110    0101001010010111    0101001010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21140 - 21144

  --0101001010011001    0101001010011010    0101001010011011    0101001010011100    0101001010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21145 - 21149

  --0101001010011110    0101001010011111    0101001010100000    0101001010100001    0101001010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21150 - 21154

  --0101001010100011    0101001010100100    0101001010100101    0101001010100110    0101001010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21155 - 21159

  --0101001010101000    0101001010101001    0101001010101010    0101001010101011    0101001010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21160 - 21164

  --0101001010101101    0101001010101110    0101001010101111    0101001010110000    0101001010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21165 - 21169

  --0101001010110010    0101001010110011    0101001010110100    0101001010110101    0101001010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21170 - 21174

  --0101001010110111    0101001010111000    0101001010111001    0101001010111010    0101001010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21175 - 21179

  --0101001010111100    0101001010111101    0101001010111110    0101001010111111    0101001011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21180 - 21184

  --0101001011000001    0101001011000010    0101001011000011    0101001011000100    0101001011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21185 - 21189

  --0101001011000110    0101001011000111    0101001011001000    0101001011001001    0101001011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21190 - 21194

  --0101001011001011    0101001011001100    0101001011001101    0101001011001110    0101001011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21195 - 21199

  --0101001011010000    0101001011010001    0101001011010010    0101001011010011    0101001011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21200 - 21204

  --0101001011010101    0101001011010110    0101001011010111    0101001011011000    0101001011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21205 - 21209

  --0101001011011010    0101001011011011    0101001011011100    0101001011011101    0101001011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21210 - 21214

  --0101001011011111    0101001011100000    0101001011100001    0101001011100010    0101001011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21215 - 21219

  --0101001011100100    0101001011100101    0101001011100110    0101001011100111    0101001011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21220 - 21224

  --0101001011101001    0101001011101010    0101001011101011    0101001011101100    0101001011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21225 - 21229

  --0101001011101110    0101001011101111    0101001011110000    0101001011110001    0101001011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21230 - 21234

  --0101001011110011    0101001011110100    0101001011110101    0101001011110110    0101001011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21235 - 21239

  --0101001011111000    0101001011111001    0101001011111010    0101001011111011    0101001011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21240 - 21244

  --0101001011111101    0101001011111110    0101001011111111    0101001100000000    0101001100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21245 - 21249

  --0101001100000010    0101001100000011    0101001100000100    0101001100000101    0101001100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21250 - 21254

  --0101001100000111    0101001100001000    0101001100001001    0101001100001010    0101001100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21255 - 21259

  --0101001100001100    0101001100001101    0101001100001110    0101001100001111    0101001100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21260 - 21264

  --0101001100010001    0101001100010010    0101001100010011    0101001100010100    0101001100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21265 - 21269

  --0101001100010110    0101001100010111    0101001100011000    0101001100011001    0101001100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21270 - 21274

  --0101001100011011    0101001100011100    0101001100011101    0101001100011110    0101001100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21275 - 21279

  --0101001100100000    0101001100100001    0101001100100010    0101001100100011    0101001100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21280 - 21284

  --0101001100100101    0101001100100110    0101001100100111    0101001100101000    0101001100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21285 - 21289

  --0101001100101010    0101001100101011    0101001100101100    0101001100101101    0101001100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21290 - 21294

  --0101001100101111    0101001100110000    0101001100110001    0101001100110010    0101001100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21295 - 21299

  --0101001100110100    0101001100110101    0101001100110110    0101001100110111    0101001100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21300 - 21304

  --0101001100111001    0101001100111010    0101001100111011    0101001100111100    0101001100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21305 - 21309

  --0101001100111110    0101001100111111    0101001101000000    0101001101000001    0101001101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21310 - 21314

  --0101001101000011    0101001101000100    0101001101000101    0101001101000110    0101001101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21315 - 21319

  --0101001101001000    0101001101001001    0101001101001010    0101001101001011    0101001101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21320 - 21324

  --0101001101001101    0101001101001110    0101001101001111    0101001101010000    0101001101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21325 - 21329

  --0101001101010010    0101001101010011    0101001101010100    0101001101010101    0101001101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21330 - 21334

  --0101001101010111    0101001101011000    0101001101011001    0101001101011010    0101001101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21335 - 21339

  --0101001101011100    0101001101011101    0101001101011110    0101001101011111    0101001101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21340 - 21344

  --0101001101100001    0101001101100010    0101001101100011    0101001101100100    0101001101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21345 - 21349

  --0101001101100110    0101001101100111    0101001101101000    0101001101101001    0101001101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21350 - 21354

  --0101001101101011    0101001101101100    0101001101101101    0101001101101110    0101001101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21355 - 21359

  --0101001101110000    0101001101110001    0101001101110010    0101001101110011    0101001101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21360 - 21364

  --0101001101110101    0101001101110110    0101001101110111    0101001101111000    0101001101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21365 - 21369

  --0101001101111010    0101001101111011    0101001101111100    0101001101111101    0101001101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21370 - 21374

  --0101001101111111    0101001110000000    0101001110000001    0101001110000010    0101001110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21375 - 21379

  --0101001110000100    0101001110000101    0101001110000110    0101001110000111    0101001110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21380 - 21384

  --0101001110001001    0101001110001010    0101001110001011    0101001110001100    0101001110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21385 - 21389

  --0101001110001110    0101001110001111    0101001110010000    0101001110010001    0101001110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21390 - 21394

  --0101001110010011    0101001110010100    0101001110010101    0101001110010110    0101001110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21395 - 21399

  --0101001110011000    0101001110011001    0101001110011010    0101001110011011    0101001110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21400 - 21404

  --0101001110011101    0101001110011110    0101001110011111    0101001110100000    0101001110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21405 - 21409

  --0101001110100010    0101001110100011    0101001110100100    0101001110100101    0101001110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21410 - 21414

  --0101001110100111    0101001110101000    0101001110101001    0101001110101010    0101001110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21415 - 21419

  --0101001110101100    0101001110101101    0101001110101110    0101001110101111    0101001110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21420 - 21424

  --0101001110110001    0101001110110010    0101001110110011    0101001110110100    0101001110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21425 - 21429

  --0101001110110110    0101001110110111    0101001110111000    0101001110111001    0101001110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21430 - 21434

  --0101001110111011    0101001110111100    0101001110111101    0101001110111110    0101001110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21435 - 21439

  --0101001111000000    0101001111000001    0101001111000010    0101001111000011    0101001111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21440 - 21444

  --0101001111000101    0101001111000110    0101001111000111    0101001111001000    0101001111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21445 - 21449

  --0101001111001010    0101001111001011    0101001111001100    0101001111001101    0101001111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21450 - 21454

  --0101001111001111    0101001111010000    0101001111010001    0101001111010010    0101001111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21455 - 21459

  --0101001111010100    0101001111010101    0101001111010110    0101001111010111    0101001111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21460 - 21464

  --0101001111011001    0101001111011010    0101001111011011    0101001111011100    0101001111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21465 - 21469

  --0101001111011110    0101001111011111    0101001111100000    0101001111100001    0101001111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21470 - 21474

  --0101001111100011    0101001111100100    0101001111100101    0101001111100110    0101001111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21475 - 21479

  --0101001111101000    0101001111101001    0101001111101010    0101001111101011    0101001111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21480 - 21484

  --0101001111101101    0101001111101110    0101001111101111    0101001111110000    0101001111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21485 - 21489

  --0101001111110010    0101001111110011    0101001111110100    0101001111110101    0101001111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21490 - 21494

  --0101001111110111    0101001111111000    0101001111111001    0101001111111010    0101001111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21495 - 21499

  --0101001111111100    0101001111111101    0101001111111110    0101001111111111    0101010000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21500 - 21504

  --0101010000000001    0101010000000010    0101010000000011    0101010000000100    0101010000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21505 - 21509

  --0101010000000110    0101010000000111    0101010000001000    0101010000001001    0101010000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21510 - 21514

  --0101010000001011    0101010000001100    0101010000001101    0101010000001110    0101010000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21515 - 21519

  --0101010000010000    0101010000010001    0101010000010010    0101010000010011    0101010000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21520 - 21524

  --0101010000010101    0101010000010110    0101010000010111    0101010000011000    0101010000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21525 - 21529

  --0101010000011010    0101010000011011    0101010000011100    0101010000011101    0101010000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21530 - 21534

  --0101010000011111    0101010000100000    0101010000100001    0101010000100010    0101010000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21535 - 21539

  --0101010000100100    0101010000100101    0101010000100110    0101010000100111    0101010000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21540 - 21544

  --0101010000101001    0101010000101010    0101010000101011    0101010000101100    0101010000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21545 - 21549

  --0101010000101110    0101010000101111    0101010000110000    0101010000110001    0101010000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21550 - 21554

  --0101010000110011    0101010000110100    0101010000110101    0101010000110110    0101010000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21555 - 21559

  --0101010000111000    0101010000111001    0101010000111010    0101010000111011    0101010000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21560 - 21564

  --0101010000111101    0101010000111110    0101010000111111    0101010001000000    0101010001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21565 - 21569

  --0101010001000010    0101010001000011    0101010001000100    0101010001000101    0101010001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21570 - 21574

  --0101010001000111    0101010001001000    0101010001001001    0101010001001010    0101010001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21575 - 21579

  --0101010001001100    0101010001001101    0101010001001110    0101010001001111    0101010001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21580 - 21584

  --0101010001010001    0101010001010010    0101010001010011    0101010001010100    0101010001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21585 - 21589

  --0101010001010110    0101010001010111    0101010001011000    0101010001011001    0101010001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21590 - 21594

  --0101010001011011    0101010001011100    0101010001011101    0101010001011110    0101010001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21595 - 21599

  --0101010001100000    0101010001100001    0101010001100010    0101010001100011    0101010001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21600 - 21604

  --0101010001100101    0101010001100110    0101010001100111    0101010001101000    0101010001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21605 - 21609

  --0101010001101010    0101010001101011    0101010001101100    0101010001101101    0101010001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21610 - 21614

  --0101010001101111    0101010001110000    0101010001110001    0101010001110010    0101010001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21615 - 21619

  --0101010001110100    0101010001110101    0101010001110110    0101010001110111    0101010001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21620 - 21624

  --0101010001111001    0101010001111010    0101010001111011    0101010001111100    0101010001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21625 - 21629

  --0101010001111110    0101010001111111    0101010010000000    0101010010000001    0101010010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21630 - 21634

  --0101010010000011    0101010010000100    0101010010000101    0101010010000110    0101010010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21635 - 21639

  --0101010010001000    0101010010001001    0101010010001010    0101010010001011    0101010010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21640 - 21644

  --0101010010001101    0101010010001110    0101010010001111    0101010010010000    0101010010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21645 - 21649

  --0101010010010010    0101010010010011    0101010010010100    0101010010010101    0101010010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21650 - 21654

  --0101010010010111    0101010010011000    0101010010011001    0101010010011010    0101010010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21655 - 21659

  --0101010010011100    0101010010011101    0101010010011110    0101010010011111    0101010010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21660 - 21664

  --0101010010100001    0101010010100010    0101010010100011    0101010010100100    0101010010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21665 - 21669

  --0101010010100110    0101010010100111    0101010010101000    0101010010101001    0101010010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21670 - 21674

  --0101010010101011    0101010010101100    0101010010101101    0101010010101110    0101010010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21675 - 21679

  --0101010010110000    0101010010110001    0101010010110010    0101010010110011    0101010010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21680 - 21684

  --0101010010110101    0101010010110110    0101010010110111    0101010010111000    0101010010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21685 - 21689

  --0101010010111010    0101010010111011    0101010010111100    0101010010111101    0101010010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21690 - 21694

  --0101010010111111    0101010011000000    0101010011000001    0101010011000010    0101010011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21695 - 21699

  --0101010011000100    0101010011000101    0101010011000110    0101010011000111    0101010011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21700 - 21704

  --0101010011001001    0101010011001010    0101010011001011    0101010011001100    0101010011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21705 - 21709

  --0101010011001110    0101010011001111    0101010011010000    0101010011010001    0101010011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21710 - 21714

  --0101010011010011    0101010011010100    0101010011010101    0101010011010110    0101010011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21715 - 21719

  --0101010011011000    0101010011011001    0101010011011010    0101010011011011    0101010011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21720 - 21724

  --0101010011011101    0101010011011110    0101010011011111    0101010011100000    0101010011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21725 - 21729

  --0101010011100010    0101010011100011    0101010011100100    0101010011100101    0101010011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21730 - 21734

  --0101010011100111    0101010011101000    0101010011101001    0101010011101010    0101010011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21735 - 21739

  --0101010011101100    0101010011101101    0101010011101110    0101010011101111    0101010011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21740 - 21744

  --0101010011110001    0101010011110010    0101010011110011    0101010011110100    0101010011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21745 - 21749

  --0101010011110110    0101010011110111    0101010011111000    0101010011111001    0101010011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21750 - 21754

  --0101010011111011    0101010011111100    0101010011111101    0101010011111110    0101010011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21755 - 21759

  --0101010100000000    0101010100000001    0101010100000010    0101010100000011    0101010100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21760 - 21764

  --0101010100000101    0101010100000110    0101010100000111    0101010100001000    0101010100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21765 - 21769

  --0101010100001010    0101010100001011    0101010100001100    0101010100001101    0101010100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21770 - 21774

  --0101010100001111    0101010100010000    0101010100010001    0101010100010010    0101010100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21775 - 21779

  --0101010100010100    0101010100010101    0101010100010110    0101010100010111    0101010100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21780 - 21784

  --0101010100011001    0101010100011010    0101010100011011    0101010100011100    0101010100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21785 - 21789

  --0101010100011110    0101010100011111    0101010100100000    0101010100100001    0101010100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21790 - 21794

  --0101010100100011    0101010100100100    0101010100100101    0101010100100110    0101010100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21795 - 21799

  --0101010100101000    0101010100101001    0101010100101010    0101010100101011    0101010100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21800 - 21804

  --0101010100101101    0101010100101110    0101010100101111    0101010100110000    0101010100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21805 - 21809

  --0101010100110010    0101010100110011    0101010100110100    0101010100110101    0101010100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21810 - 21814

  --0101010100110111    0101010100111000    0101010100111001    0101010100111010    0101010100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21815 - 21819

  --0101010100111100    0101010100111101    0101010100111110    0101010100111111    0101010101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21820 - 21824

  --0101010101000001    0101010101000010    0101010101000011    0101010101000100    0101010101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21825 - 21829

  --0101010101000110    0101010101000111    0101010101001000    0101010101001001    0101010101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21830 - 21834

  --0101010101001011    0101010101001100    0101010101001101    0101010101001110    0101010101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21835 - 21839

  --0101010101010000    0101010101010001    0101010101010010    0101010101010011    0101010101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21840 - 21844

  --0101010101010101    0101010101010110    0101010101010111    0101010101011000    0101010101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21845 - 21849

  --0101010101011010    0101010101011011    0101010101011100    0101010101011101    0101010101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21850 - 21854

  --0101010101011111    0101010101100000    0101010101100001    0101010101100010    0101010101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21855 - 21859

  --0101010101100100    0101010101100101    0101010101100110    0101010101100111    0101010101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21860 - 21864

  --0101010101101001    0101010101101010    0101010101101011    0101010101101100    0101010101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21865 - 21869

  --0101010101101110    0101010101101111    0101010101110000    0101010101110001    0101010101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21870 - 21874

  --0101010101110011    0101010101110100    0101010101110101    0101010101110110    0101010101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21875 - 21879

  --0101010101111000    0101010101111001    0101010101111010    0101010101111011    0101010101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21880 - 21884

  --0101010101111101    0101010101111110    0101010101111111    0101010110000000    0101010110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21885 - 21889

  --0101010110000010    0101010110000011    0101010110000100    0101010110000101    0101010110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21890 - 21894

  --0101010110000111    0101010110001000    0101010110001001    0101010110001010    0101010110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21895 - 21899

  --0101010110001100    0101010110001101    0101010110001110    0101010110001111    0101010110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21900 - 21904

  --0101010110010001    0101010110010010    0101010110010011    0101010110010100    0101010110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21905 - 21909

  --0101010110010110    0101010110010111    0101010110011000    0101010110011001    0101010110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21910 - 21914

  --0101010110011011    0101010110011100    0101010110011101    0101010110011110    0101010110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21915 - 21919

  --0101010110100000    0101010110100001    0101010110100010    0101010110100011    0101010110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21920 - 21924

  --0101010110100101    0101010110100110    0101010110100111    0101010110101000    0101010110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21925 - 21929

  --0101010110101010    0101010110101011    0101010110101100    0101010110101101    0101010110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21930 - 21934

  --0101010110101111    0101010110110000    0101010110110001    0101010110110010    0101010110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21935 - 21939

  --0101010110110100    0101010110110101    0101010110110110    0101010110110111    0101010110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21940 - 21944

  --0101010110111001    0101010110111010    0101010110111011    0101010110111100    0101010110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21945 - 21949

  --0101010110111110    0101010110111111    0101010111000000    0101010111000001    0101010111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21950 - 21954

  --0101010111000011    0101010111000100    0101010111000101    0101010111000110    0101010111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21955 - 21959

  --0101010111001000    0101010111001001    0101010111001010    0101010111001011    0101010111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21960 - 21964

  --0101010111001101    0101010111001110    0101010111001111    0101010111010000    0101010111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21965 - 21969

  --0101010111010010    0101010111010011    0101010111010100    0101010111010101    0101010111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21970 - 21974

  --0101010111010111    0101010111011000    0101010111011001    0101010111011010    0101010111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21975 - 21979

  --0101010111011100    0101010111011101    0101010111011110    0101010111011111    0101010111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21980 - 21984

  --0101010111100001    0101010111100010    0101010111100011    0101010111100100    0101010111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21985 - 21989

  --0101010111100110    0101010111100111    0101010111101000    0101010111101001    0101010111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21990 - 21994

  --0101010111101011    0101010111101100    0101010111101101    0101010111101110    0101010111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 21995 - 21999

  --0101010111110000    0101010111110001    0101010111110010    0101010111110011    0101010111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22000 - 22004

  --0101010111110101    0101010111110110    0101010111110111    0101010111111000    0101010111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22005 - 22009

  --0101010111111010    0101010111111011    0101010111111100    0101010111111101    0101010111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22010 - 22014

  --0101010111111111    0101011000000000    0101011000000001    0101011000000010    0101011000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22015 - 22019

  --0101011000000100    0101011000000101    0101011000000110    0101011000000111    0101011000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22020 - 22024

  --0101011000001001    0101011000001010    0101011000001011    0101011000001100    0101011000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22025 - 22029

  --0101011000001110    0101011000001111    0101011000010000    0101011000010001    0101011000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22030 - 22034

  --0101011000010011    0101011000010100    0101011000010101    0101011000010110    0101011000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22035 - 22039

  --0101011000011000    0101011000011001    0101011000011010    0101011000011011    0101011000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22040 - 22044

  --0101011000011101    0101011000011110    0101011000011111    0101011000100000    0101011000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22045 - 22049

  --0101011000100010    0101011000100011    0101011000100100    0101011000100101    0101011000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22050 - 22054

  --0101011000100111    0101011000101000    0101011000101001    0101011000101010    0101011000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22055 - 22059

  --0101011000101100    0101011000101101    0101011000101110    0101011000101111    0101011000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22060 - 22064

  --0101011000110001    0101011000110010    0101011000110011    0101011000110100    0101011000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22065 - 22069

  --0101011000110110    0101011000110111    0101011000111000    0101011000111001    0101011000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22070 - 22074

  --0101011000111011    0101011000111100    0101011000111101    0101011000111110    0101011000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22075 - 22079

  --0101011001000000    0101011001000001    0101011001000010    0101011001000011    0101011001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22080 - 22084

  --0101011001000101    0101011001000110    0101011001000111    0101011001001000    0101011001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22085 - 22089

  --0101011001001010    0101011001001011    0101011001001100    0101011001001101    0101011001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22090 - 22094

  --0101011001001111    0101011001010000    0101011001010001    0101011001010010    0101011001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22095 - 22099

  --0101011001010100    0101011001010101    0101011001010110    0101011001010111    0101011001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22100 - 22104

  --0101011001011001    0101011001011010    0101011001011011    0101011001011100    0101011001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22105 - 22109

  --0101011001011110    0101011001011111    0101011001100000    0101011001100001    0101011001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22110 - 22114

  --0101011001100011    0101011001100100    0101011001100101    0101011001100110    0101011001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22115 - 22119

  --0101011001101000    0101011001101001    0101011001101010    0101011001101011    0101011001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22120 - 22124

  --0101011001101101    0101011001101110    0101011001101111    0101011001110000    0101011001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22125 - 22129

  --0101011001110010    0101011001110011    0101011001110100    0101011001110101    0101011001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22130 - 22134

  --0101011001110111    0101011001111000    0101011001111001    0101011001111010    0101011001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22135 - 22139

  --0101011001111100    0101011001111101    0101011001111110    0101011001111111    0101011010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22140 - 22144

  --0101011010000001    0101011010000010    0101011010000011    0101011010000100    0101011010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22145 - 22149

  --0101011010000110    0101011010000111    0101011010001000    0101011010001001    0101011010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22150 - 22154

  --0101011010001011    0101011010001100    0101011010001101    0101011010001110    0101011010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22155 - 22159

  --0101011010010000    0101011010010001    0101011010010010    0101011010010011    0101011010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22160 - 22164

  --0101011010010101    0101011010010110    0101011010010111    0101011010011000    0101011010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22165 - 22169

  --0101011010011010    0101011010011011    0101011010011100    0101011010011101    0101011010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22170 - 22174

  --0101011010011111    0101011010100000    0101011010100001    0101011010100010    0101011010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22175 - 22179

  --0101011010100100    0101011010100101    0101011010100110    0101011010100111    0101011010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22180 - 22184

  --0101011010101001    0101011010101010    0101011010101011    0101011010101100    0101011010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22185 - 22189

  --0101011010101110    0101011010101111    0101011010110000    0101011010110001    0101011010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22190 - 22194

  --0101011010110011    0101011010110100    0101011010110101    0101011010110110    0101011010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22195 - 22199

  --0101011010111000    0101011010111001    0101011010111010    0101011010111011    0101011010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22200 - 22204

  --0101011010111101    0101011010111110    0101011010111111    0101011011000000    0101011011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22205 - 22209

  --0101011011000010    0101011011000011    0101011011000100    0101011011000101    0101011011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22210 - 22214

  --0101011011000111    0101011011001000    0101011011001001    0101011011001010    0101011011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22215 - 22219

  --0101011011001100    0101011011001101    0101011011001110    0101011011001111    0101011011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22220 - 22224

  --0101011011010001    0101011011010010    0101011011010011    0101011011010100    0101011011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22225 - 22229

  --0101011011010110    0101011011010111    0101011011011000    0101011011011001    0101011011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22230 - 22234

  --0101011011011011    0101011011011100    0101011011011101    0101011011011110    0101011011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22235 - 22239

  --0101011011100000    0101011011100001    0101011011100010    0101011011100011    0101011011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22240 - 22244

  --0101011011100101    0101011011100110    0101011011100111    0101011011101000    0101011011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22245 - 22249

  --0101011011101010    0101011011101011    0101011011101100    0101011011101101    0101011011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22250 - 22254

  --0101011011101111    0101011011110000    0101011011110001    0101011011110010    0101011011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22255 - 22259

  --0101011011110100    0101011011110101    0101011011110110    0101011011110111    0101011011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22260 - 22264

  --0101011011111001    0101011011111010    0101011011111011    0101011011111100    0101011011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22265 - 22269

  --0101011011111110    0101011011111111    0101011100000000    0101011100000001    0101011100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22270 - 22274

  --0101011100000011    0101011100000100    0101011100000101    0101011100000110    0101011100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22275 - 22279

  --0101011100001000    0101011100001001    0101011100001010    0101011100001011    0101011100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22280 - 22284

  --0101011100001101    0101011100001110    0101011100001111    0101011100010000    0101011100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22285 - 22289

  --0101011100010010    0101011100010011    0101011100010100    0101011100010101    0101011100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22290 - 22294

  --0101011100010111    0101011100011000    0101011100011001    0101011100011010    0101011100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22295 - 22299

  --0101011100011100    0101011100011101    0101011100011110    0101011100011111    0101011100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22300 - 22304

  --0101011100100001    0101011100100010    0101011100100011    0101011100100100    0101011100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22305 - 22309

  --0101011100100110    0101011100100111    0101011100101000    0101011100101001    0101011100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22310 - 22314

  --0101011100101011    0101011100101100    0101011100101101    0101011100101110    0101011100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22315 - 22319

  --0101011100110000    0101011100110001    0101011100110010    0101011100110011    0101011100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22320 - 22324

  --0101011100110101    0101011100110110    0101011100110111    0101011100111000    0101011100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22325 - 22329

  --0101011100111010    0101011100111011    0101011100111100    0101011100111101    0101011100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22330 - 22334

  --0101011100111111    0101011101000000    0101011101000001    0101011101000010    0101011101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22335 - 22339

  --0101011101000100    0101011101000101    0101011101000110    0101011101000111    0101011101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22340 - 22344

  --0101011101001001    0101011101001010    0101011101001011    0101011101001100    0101011101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22345 - 22349

  --0101011101001110    0101011101001111    0101011101010000    0101011101010001    0101011101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22350 - 22354

  --0101011101010011    0101011101010100    0101011101010101    0101011101010110    0101011101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22355 - 22359

  --0101011101011000    0101011101011001    0101011101011010    0101011101011011    0101011101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22360 - 22364

  --0101011101011101    0101011101011110    0101011101011111    0101011101100000    0101011101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22365 - 22369

  --0101011101100010    0101011101100011    0101011101100100    0101011101100101    0101011101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22370 - 22374

  --0101011101100111    0101011101101000    0101011101101001    0101011101101010    0101011101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22375 - 22379

  --0101011101101100    0101011101101101    0101011101101110    0101011101101111    0101011101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22380 - 22384

  --0101011101110001    0101011101110010    0101011101110011    0101011101110100    0101011101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22385 - 22389

  --0101011101110110    0101011101110111    0101011101111000    0101011101111001    0101011101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22390 - 22394

  --0101011101111011    0101011101111100    0101011101111101    0101011101111110    0101011101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22395 - 22399

  --0101011110000000    0101011110000001    0101011110000010    0101011110000011    0101011110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22400 - 22404

  --0101011110000101    0101011110000110    0101011110000111    0101011110001000    0101011110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22405 - 22409

  --0101011110001010    0101011110001011    0101011110001100    0101011110001101    0101011110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22410 - 22414

  --0101011110001111    0101011110010000    0101011110010001    0101011110010010    0101011110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22415 - 22419

  --0101011110010100    0101011110010101    0101011110010110    0101011110010111    0101011110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22420 - 22424

  --0101011110011001    0101011110011010    0101011110011011    0101011110011100    0101011110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22425 - 22429

  --0101011110011110    0101011110011111    0101011110100000    0101011110100001    0101011110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22430 - 22434

  --0101011110100011    0101011110100100    0101011110100101    0101011110100110    0101011110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22435 - 22439

  --0101011110101000    0101011110101001    0101011110101010    0101011110101011    0101011110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22440 - 22444

  --0101011110101101    0101011110101110    0101011110101111    0101011110110000    0101011110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22445 - 22449

  --0101011110110010    0101011110110011    0101011110110100    0101011110110101    0101011110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22450 - 22454

  --0101011110110111    0101011110111000    0101011110111001    0101011110111010    0101011110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22455 - 22459

  --0101011110111100    0101011110111101    0101011110111110    0101011110111111    0101011111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22460 - 22464

  --0101011111000001    0101011111000010    0101011111000011    0101011111000100    0101011111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22465 - 22469

  --0101011111000110    0101011111000111    0101011111001000    0101011111001001    0101011111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22470 - 22474

  --0101011111001011    0101011111001100    0101011111001101    0101011111001110    0101011111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22475 - 22479

  --0101011111010000    0101011111010001    0101011111010010    0101011111010011    0101011111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22480 - 22484

  --0101011111010101    0101011111010110    0101011111010111    0101011111011000    0101011111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22485 - 22489

  --0101011111011010    0101011111011011    0101011111011100    0101011111011101    0101011111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22490 - 22494

  --0101011111011111    0101011111100000    0101011111100001    0101011111100010    0101011111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22495 - 22499

  --0101011111100100    0101011111100101    0101011111100110    0101011111100111    0101011111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22500 - 22504

  --0101011111101001    0101011111101010    0101011111101011    0101011111101100    0101011111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22505 - 22509

  --0101011111101110    0101011111101111    0101011111110000    0101011111110001    0101011111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22510 - 22514

  --0101011111110011    0101011111110100    0101011111110101    0101011111110110    0101011111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22515 - 22519

  --0101011111111000    0101011111111001    0101011111111010    0101011111111011    0101011111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22520 - 22524

  --0101011111111101    0101011111111110    0101011111111111    0101100000000000    0101100000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22525 - 22529

  --0101100000000010    0101100000000011    0101100000000100    0101100000000101    0101100000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22530 - 22534

  --0101100000000111    0101100000001000    0101100000001001    0101100000001010    0101100000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22535 - 22539

  --0101100000001100    0101100000001101    0101100000001110    0101100000001111    0101100000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22540 - 22544

  --0101100000010001    0101100000010010    0101100000010011    0101100000010100    0101100000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22545 - 22549

  --0101100000010110    0101100000010111    0101100000011000    0101100000011001    0101100000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22550 - 22554

  --0101100000011011    0101100000011100    0101100000011101    0101100000011110    0101100000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22555 - 22559

  --0101100000100000    0101100000100001    0101100000100010    0101100000100011    0101100000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22560 - 22564

  --0101100000100101    0101100000100110    0101100000100111    0101100000101000    0101100000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22565 - 22569

  --0101100000101010    0101100000101011    0101100000101100    0101100000101101    0101100000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22570 - 22574

  --0101100000101111    0101100000110000    0101100000110001    0101100000110010    0101100000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22575 - 22579

  --0101100000110100    0101100000110101    0101100000110110    0101100000110111    0101100000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22580 - 22584

  --0101100000111001    0101100000111010    0101100000111011    0101100000111100    0101100000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22585 - 22589

  --0101100000111110    0101100000111111    0101100001000000    0101100001000001    0101100001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22590 - 22594

  --0101100001000011    0101100001000100    0101100001000101    0101100001000110    0101100001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22595 - 22599

  --0101100001001000    0101100001001001    0101100001001010    0101100001001011    0101100001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22600 - 22604

  --0101100001001101    0101100001001110    0101100001001111    0101100001010000    0101100001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22605 - 22609

  --0101100001010010    0101100001010011    0101100001010100    0101100001010101    0101100001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22610 - 22614

  --0101100001010111    0101100001011000    0101100001011001    0101100001011010    0101100001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22615 - 22619

  --0101100001011100    0101100001011101    0101100001011110    0101100001011111    0101100001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22620 - 22624

  --0101100001100001    0101100001100010    0101100001100011    0101100001100100    0101100001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22625 - 22629

  --0101100001100110    0101100001100111    0101100001101000    0101100001101001    0101100001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22630 - 22634

  --0101100001101011    0101100001101100    0101100001101101    0101100001101110    0101100001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22635 - 22639

  --0101100001110000    0101100001110001    0101100001110010    0101100001110011    0101100001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22640 - 22644

  --0101100001110101    0101100001110110    0101100001110111    0101100001111000    0101100001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22645 - 22649

  --0101100001111010    0101100001111011    0101100001111100    0101100001111101    0101100001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22650 - 22654

  --0101100001111111    0101100010000000    0101100010000001    0101100010000010    0101100010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22655 - 22659

  --0101100010000100    0101100010000101    0101100010000110    0101100010000111    0101100010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22660 - 22664

  --0101100010001001    0101100010001010    0101100010001011    0101100010001100    0101100010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22665 - 22669

  --0101100010001110    0101100010001111    0101100010010000    0101100010010001    0101100010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22670 - 22674

  --0101100010010011    0101100010010100    0101100010010101    0101100010010110    0101100010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22675 - 22679

  --0101100010011000    0101100010011001    0101100010011010    0101100010011011    0101100010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22680 - 22684

  --0101100010011101    0101100010011110    0101100010011111    0101100010100000    0101100010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22685 - 22689

  --0101100010100010    0101100010100011    0101100010100100    0101100010100101    0101100010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22690 - 22694

  --0101100010100111    0101100010101000    0101100010101001    0101100010101010    0101100010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22695 - 22699

  --0101100010101100    0101100010101101    0101100010101110    0101100010101111    0101100010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22700 - 22704

  --0101100010110001    0101100010110010    0101100010110011    0101100010110100    0101100010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22705 - 22709

  --0101100010110110    0101100010110111    0101100010111000    0101100010111001    0101100010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22710 - 22714

  --0101100010111011    0101100010111100    0101100010111101    0101100010111110    0101100010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22715 - 22719

  --0101100011000000    0101100011000001    0101100011000010    0101100011000011    0101100011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22720 - 22724

  --0101100011000101    0101100011000110    0101100011000111    0101100011001000    0101100011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22725 - 22729

  --0101100011001010    0101100011001011    0101100011001100    0101100011001101    0101100011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22730 - 22734

  --0101100011001111    0101100011010000    0101100011010001    0101100011010010    0101100011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22735 - 22739

  --0101100011010100    0101100011010101    0101100011010110    0101100011010111    0101100011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22740 - 22744

  --0101100011011001    0101100011011010    0101100011011011    0101100011011100    0101100011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22745 - 22749

  --0101100011011110    0101100011011111    0101100011100000    0101100011100001    0101100011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22750 - 22754

  --0101100011100011    0101100011100100    0101100011100101    0101100011100110    0101100011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22755 - 22759

  --0101100011101000    0101100011101001    0101100011101010    0101100011101011    0101100011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22760 - 22764

  --0101100011101101    0101100011101110    0101100011101111    0101100011110000    0101100011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22765 - 22769

  --0101100011110010    0101100011110011    0101100011110100    0101100011110101    0101100011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22770 - 22774

  --0101100011110111    0101100011111000    0101100011111001    0101100011111010    0101100011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22775 - 22779

  --0101100011111100    0101100011111101    0101100011111110    0101100011111111    0101100100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22780 - 22784

  --0101100100000001    0101100100000010    0101100100000011    0101100100000100    0101100100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22785 - 22789

  --0101100100000110    0101100100000111    0101100100001000    0101100100001001    0101100100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22790 - 22794

  --0101100100001011    0101100100001100    0101100100001101    0101100100001110    0101100100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22795 - 22799

  --0101100100010000    0101100100010001    0101100100010010    0101100100010011    0101100100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22800 - 22804

  --0101100100010101    0101100100010110    0101100100010111    0101100100011000    0101100100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22805 - 22809

  --0101100100011010    0101100100011011    0101100100011100    0101100100011101    0101100100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22810 - 22814

  --0101100100011111    0101100100100000    0101100100100001    0101100100100010    0101100100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22815 - 22819

  --0101100100100100    0101100100100101    0101100100100110    0101100100100111    0101100100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22820 - 22824

  --0101100100101001    0101100100101010    0101100100101011    0101100100101100    0101100100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22825 - 22829

  --0101100100101110    0101100100101111    0101100100110000    0101100100110001    0101100100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22830 - 22834

  --0101100100110011    0101100100110100    0101100100110101    0101100100110110    0101100100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22835 - 22839

  --0101100100111000    0101100100111001    0101100100111010    0101100100111011    0101100100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22840 - 22844

  --0101100100111101    0101100100111110    0101100100111111    0101100101000000    0101100101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22845 - 22849

  --0101100101000010    0101100101000011    0101100101000100    0101100101000101    0101100101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22850 - 22854

  --0101100101000111    0101100101001000    0101100101001001    0101100101001010    0101100101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22855 - 22859

  --0101100101001100    0101100101001101    0101100101001110    0101100101001111    0101100101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22860 - 22864

  --0101100101010001    0101100101010010    0101100101010011    0101100101010100    0101100101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22865 - 22869

  --0101100101010110    0101100101010111    0101100101011000    0101100101011001    0101100101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22870 - 22874

  --0101100101011011    0101100101011100    0101100101011101    0101100101011110    0101100101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22875 - 22879

  --0101100101100000    0101100101100001    0101100101100010    0101100101100011    0101100101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22880 - 22884

  --0101100101100101    0101100101100110    0101100101100111    0101100101101000    0101100101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22885 - 22889

  --0101100101101010    0101100101101011    0101100101101100    0101100101101101    0101100101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22890 - 22894

  --0101100101101111    0101100101110000    0101100101110001    0101100101110010    0101100101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22895 - 22899

  --0101100101110100    0101100101110101    0101100101110110    0101100101110111    0101100101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22900 - 22904

  --0101100101111001    0101100101111010    0101100101111011    0101100101111100    0101100101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22905 - 22909

  --0101100101111110    0101100101111111    0101100110000000    0101100110000001    0101100110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22910 - 22914

  --0101100110000011    0101100110000100    0101100110000101    0101100110000110    0101100110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22915 - 22919

  --0101100110001000    0101100110001001    0101100110001010    0101100110001011    0101100110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22920 - 22924

  --0101100110001101    0101100110001110    0101100110001111    0101100110010000    0101100110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22925 - 22929

  --0101100110010010    0101100110010011    0101100110010100    0101100110010101    0101100110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22930 - 22934

  --0101100110010111    0101100110011000    0101100110011001    0101100110011010    0101100110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22935 - 22939

  --0101100110011100    0101100110011101    0101100110011110    0101100110011111    0101100110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22940 - 22944

  --0101100110100001    0101100110100010    0101100110100011    0101100110100100    0101100110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22945 - 22949

  --0101100110100110    0101100110100111    0101100110101000    0101100110101001    0101100110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22950 - 22954

  --0101100110101011    0101100110101100    0101100110101101    0101100110101110    0101100110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22955 - 22959

  --0101100110110000    0101100110110001    0101100110110010    0101100110110011    0101100110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22960 - 22964

  --0101100110110101    0101100110110110    0101100110110111    0101100110111000    0101100110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22965 - 22969

  --0101100110111010    0101100110111011    0101100110111100    0101100110111101    0101100110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22970 - 22974

  --0101100110111111    0101100111000000    0101100111000001    0101100111000010    0101100111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22975 - 22979

  --0101100111000100    0101100111000101    0101100111000110    0101100111000111    0101100111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22980 - 22984

  --0101100111001001    0101100111001010    0101100111001011    0101100111001100    0101100111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22985 - 22989

  --0101100111001110    0101100111001111    0101100111010000    0101100111010001    0101100111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22990 - 22994

  --0101100111010011    0101100111010100    0101100111010101    0101100111010110    0101100111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 22995 - 22999

  --0101100111011000    0101100111011001    0101100111011010    0101100111011011    0101100111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23000 - 23004

  --0101100111011101    0101100111011110    0101100111011111    0101100111100000    0101100111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23005 - 23009

  --0101100111100010    0101100111100011    0101100111100100    0101100111100101    0101100111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23010 - 23014

  --0101100111100111    0101100111101000    0101100111101001    0101100111101010    0101100111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23015 - 23019

  --0101100111101100    0101100111101101    0101100111101110    0101100111101111    0101100111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23020 - 23024

  --0101100111110001    0101100111110010    0101100111110011    0101100111110100    0101100111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23025 - 23029

  --0101100111110110    0101100111110111    0101100111111000    0101100111111001    0101100111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23030 - 23034

  --0101100111111011    0101100111111100    0101100111111101    0101100111111110    0101100111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23035 - 23039

  --0101101000000000    0101101000000001    0101101000000010    0101101000000011    0101101000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23040 - 23044

  --0101101000000101    0101101000000110    0101101000000111    0101101000001000    0101101000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23045 - 23049

  --0101101000001010    0101101000001011    0101101000001100    0101101000001101    0101101000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23050 - 23054

  --0101101000001111    0101101000010000    0101101000010001    0101101000010010    0101101000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23055 - 23059

  --0101101000010100    0101101000010101    0101101000010110    0101101000010111    0101101000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23060 - 23064

  --0101101000011001    0101101000011010    0101101000011011    0101101000011100    0101101000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23065 - 23069

  --0101101000011110    0101101000011111    0101101000100000    0101101000100001    0101101000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23070 - 23074

  --0101101000100011    0101101000100100    0101101000100101    0101101000100110    0101101000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23075 - 23079

  --0101101000101000    0101101000101001    0101101000101010    0101101000101011    0101101000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23080 - 23084

  --0101101000101101    0101101000101110    0101101000101111    0101101000110000    0101101000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23085 - 23089

  --0101101000110010    0101101000110011    0101101000110100    0101101000110101    0101101000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23090 - 23094

  --0101101000110111    0101101000111000    0101101000111001    0101101000111010    0101101000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23095 - 23099

  --0101101000111100    0101101000111101    0101101000111110    0101101000111111    0101101001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23100 - 23104

  --0101101001000001    0101101001000010    0101101001000011    0101101001000100    0101101001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23105 - 23109

  --0101101001000110    0101101001000111    0101101001001000    0101101001001001    0101101001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23110 - 23114

  --0101101001001011    0101101001001100    0101101001001101    0101101001001110    0101101001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23115 - 23119

  --0101101001010000    0101101001010001    0101101001010010    0101101001010011    0101101001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23120 - 23124

  --0101101001010101    0101101001010110    0101101001010111    0101101001011000    0101101001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23125 - 23129

  --0101101001011010    0101101001011011    0101101001011100    0101101001011101    0101101001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23130 - 23134

  --0101101001011111    0101101001100000    0101101001100001    0101101001100010    0101101001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23135 - 23139

  --0101101001100100    0101101001100101    0101101001100110    0101101001100111    0101101001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23140 - 23144

  --0101101001101001    0101101001101010    0101101001101011    0101101001101100    0101101001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23145 - 23149

  --0101101001101110    0101101001101111    0101101001110000    0101101001110001    0101101001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23150 - 23154

  --0101101001110011    0101101001110100    0101101001110101    0101101001110110    0101101001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23155 - 23159

  --0101101001111000    0101101001111001    0101101001111010    0101101001111011    0101101001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23160 - 23164

  --0101101001111101    0101101001111110    0101101001111111    0101101010000000    0101101010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23165 - 23169

  --0101101010000010    0101101010000011    0101101010000100    0101101010000101    0101101010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23170 - 23174

  --0101101010000111    0101101010001000    0101101010001001    0101101010001010    0101101010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23175 - 23179

  --0101101010001100    0101101010001101    0101101010001110    0101101010001111    0101101010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23180 - 23184

  --0101101010010001    0101101010010010    0101101010010011    0101101010010100    0101101010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23185 - 23189

  --0101101010010110    0101101010010111    0101101010011000    0101101010011001    0101101010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23190 - 23194

  --0101101010011011    0101101010011100    0101101010011101    0101101010011110    0101101010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23195 - 23199

  --0101101010100000    0101101010100001    0101101010100010    0101101010100011    0101101010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23200 - 23204

  --0101101010100101    0101101010100110    0101101010100111    0101101010101000    0101101010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23205 - 23209

  --0101101010101010    0101101010101011    0101101010101100    0101101010101101    0101101010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23210 - 23214

  --0101101010101111    0101101010110000    0101101010110001    0101101010110010    0101101010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23215 - 23219

  --0101101010110100    0101101010110101    0101101010110110    0101101010110111    0101101010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23220 - 23224

  --0101101010111001    0101101010111010    0101101010111011    0101101010111100    0101101010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23225 - 23229

  --0101101010111110    0101101010111111    0101101011000000    0101101011000001    0101101011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23230 - 23234

  --0101101011000011    0101101011000100    0101101011000101    0101101011000110    0101101011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23235 - 23239

  --0101101011001000    0101101011001001    0101101011001010    0101101011001011    0101101011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23240 - 23244

  --0101101011001101    0101101011001110    0101101011001111    0101101011010000    0101101011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23245 - 23249

  --0101101011010010    0101101011010011    0101101011010100    0101101011010101    0101101011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23250 - 23254

  --0101101011010111    0101101011011000    0101101011011001    0101101011011010    0101101011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23255 - 23259

  --0101101011011100    0101101011011101    0101101011011110    0101101011011111    0101101011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23260 - 23264

  --0101101011100001    0101101011100010    0101101011100011    0101101011100100    0101101011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23265 - 23269

  --0101101011100110    0101101011100111    0101101011101000    0101101011101001    0101101011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23270 - 23274

  --0101101011101011    0101101011101100    0101101011101101    0101101011101110    0101101011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23275 - 23279

  --0101101011110000    0101101011110001    0101101011110010    0101101011110011    0101101011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23280 - 23284

  --0101101011110101    0101101011110110    0101101011110111    0101101011111000    0101101011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23285 - 23289

  --0101101011111010    0101101011111011    0101101011111100    0101101011111101    0101101011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23290 - 23294

  --0101101011111111    0101101100000000    0101101100000001    0101101100000010    0101101100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23295 - 23299

  --0101101100000100    0101101100000101    0101101100000110    0101101100000111    0101101100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23300 - 23304

  --0101101100001001    0101101100001010    0101101100001011    0101101100001100    0101101100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23305 - 23309

  --0101101100001110    0101101100001111    0101101100010000    0101101100010001    0101101100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23310 - 23314

  --0101101100010011    0101101100010100    0101101100010101    0101101100010110    0101101100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23315 - 23319

  --0101101100011000    0101101100011001    0101101100011010    0101101100011011    0101101100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23320 - 23324

  --0101101100011101    0101101100011110    0101101100011111    0101101100100000    0101101100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23325 - 23329

  --0101101100100010    0101101100100011    0101101100100100    0101101100100101    0101101100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23330 - 23334

  --0101101100100111    0101101100101000    0101101100101001    0101101100101010    0101101100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23335 - 23339

  --0101101100101100    0101101100101101    0101101100101110    0101101100101111    0101101100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23340 - 23344

  --0101101100110001    0101101100110010    0101101100110011    0101101100110100    0101101100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23345 - 23349

  --0101101100110110    0101101100110111    0101101100111000    0101101100111001    0101101100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23350 - 23354

  --0101101100111011    0101101100111100    0101101100111101    0101101100111110    0101101100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23355 - 23359

  --0101101101000000    0101101101000001    0101101101000010    0101101101000011    0101101101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23360 - 23364

  --0101101101000101    0101101101000110    0101101101000111    0101101101001000    0101101101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23365 - 23369

  --0101101101001010    0101101101001011    0101101101001100    0101101101001101    0101101101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23370 - 23374

  --0101101101001111    0101101101010000    0101101101010001    0101101101010010    0101101101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23375 - 23379

  --0101101101010100    0101101101010101    0101101101010110    0101101101010111    0101101101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23380 - 23384

  --0101101101011001    0101101101011010    0101101101011011    0101101101011100    0101101101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23385 - 23389

  --0101101101011110    0101101101011111    0101101101100000    0101101101100001    0101101101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23390 - 23394

  --0101101101100011    0101101101100100    0101101101100101    0101101101100110    0101101101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23395 - 23399

  --0101101101101000    0101101101101001    0101101101101010    0101101101101011    0101101101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23400 - 23404

  --0101101101101101    0101101101101110    0101101101101111    0101101101110000    0101101101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23405 - 23409

  --0101101101110010    0101101101110011    0101101101110100    0101101101110101    0101101101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23410 - 23414

  --0101101101110111    0101101101111000    0101101101111001    0101101101111010    0101101101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23415 - 23419

  --0101101101111100    0101101101111101    0101101101111110    0101101101111111    0101101110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23420 - 23424

  --0101101110000001    0101101110000010    0101101110000011    0101101110000100    0101101110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23425 - 23429

  --0101101110000110    0101101110000111    0101101110001000    0101101110001001    0101101110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23430 - 23434

  --0101101110001011    0101101110001100    0101101110001101    0101101110001110    0101101110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23435 - 23439

  --0101101110010000    0101101110010001    0101101110010010    0101101110010011    0101101110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23440 - 23444

  --0101101110010101    0101101110010110    0101101110010111    0101101110011000    0101101110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23445 - 23449

  --0101101110011010    0101101110011011    0101101110011100    0101101110011101    0101101110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23450 - 23454

  --0101101110011111    0101101110100000    0101101110100001    0101101110100010    0101101110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23455 - 23459

  --0101101110100100    0101101110100101    0101101110100110    0101101110100111    0101101110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23460 - 23464

  --0101101110101001    0101101110101010    0101101110101011    0101101110101100    0101101110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23465 - 23469

  --0101101110101110    0101101110101111    0101101110110000    0101101110110001    0101101110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23470 - 23474

  --0101101110110011    0101101110110100    0101101110110101    0101101110110110    0101101110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23475 - 23479

  --0101101110111000    0101101110111001    0101101110111010    0101101110111011    0101101110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23480 - 23484

  --0101101110111101    0101101110111110    0101101110111111    0101101111000000    0101101111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23485 - 23489

  --0101101111000010    0101101111000011    0101101111000100    0101101111000101    0101101111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23490 - 23494

  --0101101111000111    0101101111001000    0101101111001001    0101101111001010    0101101111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23495 - 23499

  --0101101111001100    0101101111001101    0101101111001110    0101101111001111    0101101111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23500 - 23504

  --0101101111010001    0101101111010010    0101101111010011    0101101111010100    0101101111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23505 - 23509

  --0101101111010110    0101101111010111    0101101111011000    0101101111011001    0101101111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23510 - 23514

  --0101101111011011    0101101111011100    0101101111011101    0101101111011110    0101101111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23515 - 23519

  --0101101111100000    0101101111100001    0101101111100010    0101101111100011    0101101111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23520 - 23524

  --0101101111100101    0101101111100110    0101101111100111    0101101111101000    0101101111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23525 - 23529

  --0101101111101010    0101101111101011    0101101111101100    0101101111101101    0101101111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23530 - 23534

  --0101101111101111    0101101111110000    0101101111110001    0101101111110010    0101101111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23535 - 23539

  --0101101111110100    0101101111110101    0101101111110110    0101101111110111    0101101111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23540 - 23544

  --0101101111111001    0101101111111010    0101101111111011    0101101111111100    0101101111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23545 - 23549

  --0101101111111110    0101101111111111    0101110000000000    0101110000000001    0101110000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23550 - 23554

  --0101110000000011    0101110000000100    0101110000000101    0101110000000110    0101110000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23555 - 23559

  --0101110000001000    0101110000001001    0101110000001010    0101110000001011    0101110000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23560 - 23564

  --0101110000001101    0101110000001110    0101110000001111    0101110000010000    0101110000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23565 - 23569

  --0101110000010010    0101110000010011    0101110000010100    0101110000010101    0101110000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23570 - 23574

  --0101110000010111    0101110000011000    0101110000011001    0101110000011010    0101110000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23575 - 23579

  --0101110000011100    0101110000011101    0101110000011110    0101110000011111    0101110000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23580 - 23584

  --0101110000100001    0101110000100010    0101110000100011    0101110000100100    0101110000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23585 - 23589

  --0101110000100110    0101110000100111    0101110000101000    0101110000101001    0101110000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23590 - 23594

  --0101110000101011    0101110000101100    0101110000101101    0101110000101110    0101110000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23595 - 23599

  --0101110000110000    0101110000110001    0101110000110010    0101110000110011    0101110000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23600 - 23604

  --0101110000110101    0101110000110110    0101110000110111    0101110000111000    0101110000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23605 - 23609

  --0101110000111010    0101110000111011    0101110000111100    0101110000111101    0101110000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23610 - 23614

  --0101110000111111    0101110001000000    0101110001000001    0101110001000010    0101110001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23615 - 23619

  --0101110001000100    0101110001000101    0101110001000110    0101110001000111    0101110001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23620 - 23624

  --0101110001001001    0101110001001010    0101110001001011    0101110001001100    0101110001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23625 - 23629

  --0101110001001110    0101110001001111    0101110001010000    0101110001010001    0101110001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23630 - 23634

  --0101110001010011    0101110001010100    0101110001010101    0101110001010110    0101110001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23635 - 23639

  --0101110001011000    0101110001011001    0101110001011010    0101110001011011    0101110001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23640 - 23644

  --0101110001011101    0101110001011110    0101110001011111    0101110001100000    0101110001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23645 - 23649

  --0101110001100010    0101110001100011    0101110001100100    0101110001100101    0101110001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23650 - 23654

  --0101110001100111    0101110001101000    0101110001101001    0101110001101010    0101110001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23655 - 23659

  --0101110001101100    0101110001101101    0101110001101110    0101110001101111    0101110001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23660 - 23664

  --0101110001110001    0101110001110010    0101110001110011    0101110001110100    0101110001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23665 - 23669

  --0101110001110110    0101110001110111    0101110001111000    0101110001111001    0101110001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23670 - 23674

  --0101110001111011    0101110001111100    0101110001111101    0101110001111110    0101110001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23675 - 23679

  --0101110010000000    0101110010000001    0101110010000010    0101110010000011    0101110010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23680 - 23684

  --0101110010000101    0101110010000110    0101110010000111    0101110010001000    0101110010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23685 - 23689

  --0101110010001010    0101110010001011    0101110010001100    0101110010001101    0101110010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23690 - 23694

  --0101110010001111    0101110010010000    0101110010010001    0101110010010010    0101110010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23695 - 23699

  --0101110010010100    0101110010010101    0101110010010110    0101110010010111    0101110010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23700 - 23704

  --0101110010011001    0101110010011010    0101110010011011    0101110010011100    0101110010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23705 - 23709

  --0101110010011110    0101110010011111    0101110010100000    0101110010100001    0101110010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23710 - 23714

  --0101110010100011    0101110010100100    0101110010100101    0101110010100110    0101110010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23715 - 23719

  --0101110010101000    0101110010101001    0101110010101010    0101110010101011    0101110010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23720 - 23724

  --0101110010101101    0101110010101110    0101110010101111    0101110010110000    0101110010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23725 - 23729

  --0101110010110010    0101110010110011    0101110010110100    0101110010110101    0101110010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23730 - 23734

  --0101110010110111    0101110010111000    0101110010111001    0101110010111010    0101110010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23735 - 23739

  --0101110010111100    0101110010111101    0101110010111110    0101110010111111    0101110011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23740 - 23744

  --0101110011000001    0101110011000010    0101110011000011    0101110011000100    0101110011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23745 - 23749

  --0101110011000110    0101110011000111    0101110011001000    0101110011001001    0101110011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23750 - 23754

  --0101110011001011    0101110011001100    0101110011001101    0101110011001110    0101110011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23755 - 23759

  --0101110011010000    0101110011010001    0101110011010010    0101110011010011    0101110011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23760 - 23764

  --0101110011010101    0101110011010110    0101110011010111    0101110011011000    0101110011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23765 - 23769

  --0101110011011010    0101110011011011    0101110011011100    0101110011011101    0101110011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23770 - 23774

  --0101110011011111    0101110011100000    0101110011100001    0101110011100010    0101110011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23775 - 23779

  --0101110011100100    0101110011100101    0101110011100110    0101110011100111    0101110011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23780 - 23784

  --0101110011101001    0101110011101010    0101110011101011    0101110011101100    0101110011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23785 - 23789

  --0101110011101110    0101110011101111    0101110011110000    0101110011110001    0101110011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23790 - 23794

  --0101110011110011    0101110011110100    0101110011110101    0101110011110110    0101110011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23795 - 23799

  --0101110011111000    0101110011111001    0101110011111010    0101110011111011    0101110011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23800 - 23804

  --0101110011111101    0101110011111110    0101110011111111    0101110100000000    0101110100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23805 - 23809

  --0101110100000010    0101110100000011    0101110100000100    0101110100000101    0101110100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23810 - 23814

  --0101110100000111    0101110100001000    0101110100001001    0101110100001010    0101110100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23815 - 23819

  --0101110100001100    0101110100001101    0101110100001110    0101110100001111    0101110100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23820 - 23824

  --0101110100010001    0101110100010010    0101110100010011    0101110100010100    0101110100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23825 - 23829

  --0101110100010110    0101110100010111    0101110100011000    0101110100011001    0101110100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23830 - 23834

  --0101110100011011    0101110100011100    0101110100011101    0101110100011110    0101110100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23835 - 23839

  --0101110100100000    0101110100100001    0101110100100010    0101110100100011    0101110100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23840 - 23844

  --0101110100100101    0101110100100110    0101110100100111    0101110100101000    0101110100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23845 - 23849

  --0101110100101010    0101110100101011    0101110100101100    0101110100101101    0101110100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23850 - 23854

  --0101110100101111    0101110100110000    0101110100110001    0101110100110010    0101110100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23855 - 23859

  --0101110100110100    0101110100110101    0101110100110110    0101110100110111    0101110100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23860 - 23864

  --0101110100111001    0101110100111010    0101110100111011    0101110100111100    0101110100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23865 - 23869

  --0101110100111110    0101110100111111    0101110101000000    0101110101000001    0101110101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23870 - 23874

  --0101110101000011    0101110101000100    0101110101000101    0101110101000110    0101110101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23875 - 23879

  --0101110101001000    0101110101001001    0101110101001010    0101110101001011    0101110101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23880 - 23884

  --0101110101001101    0101110101001110    0101110101001111    0101110101010000    0101110101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23885 - 23889

  --0101110101010010    0101110101010011    0101110101010100    0101110101010101    0101110101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23890 - 23894

  --0101110101010111    0101110101011000    0101110101011001    0101110101011010    0101110101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23895 - 23899

  --0101110101011100    0101110101011101    0101110101011110    0101110101011111    0101110101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23900 - 23904

  --0101110101100001    0101110101100010    0101110101100011    0101110101100100    0101110101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23905 - 23909

  --0101110101100110    0101110101100111    0101110101101000    0101110101101001    0101110101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23910 - 23914

  --0101110101101011    0101110101101100    0101110101101101    0101110101101110    0101110101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23915 - 23919

  --0101110101110000    0101110101110001    0101110101110010    0101110101110011    0101110101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23920 - 23924

  --0101110101110101    0101110101110110    0101110101110111    0101110101111000    0101110101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23925 - 23929

  --0101110101111010    0101110101111011    0101110101111100    0101110101111101    0101110101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23930 - 23934

  --0101110101111111    0101110110000000    0101110110000001    0101110110000010    0101110110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23935 - 23939

  --0101110110000100    0101110110000101    0101110110000110    0101110110000111    0101110110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23940 - 23944

  --0101110110001001    0101110110001010    0101110110001011    0101110110001100    0101110110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23945 - 23949

  --0101110110001110    0101110110001111    0101110110010000    0101110110010001    0101110110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23950 - 23954

  --0101110110010011    0101110110010100    0101110110010101    0101110110010110    0101110110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23955 - 23959

  --0101110110011000    0101110110011001    0101110110011010    0101110110011011    0101110110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23960 - 23964

  --0101110110011101    0101110110011110    0101110110011111    0101110110100000    0101110110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23965 - 23969

  --0101110110100010    0101110110100011    0101110110100100    0101110110100101    0101110110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23970 - 23974

  --0101110110100111    0101110110101000    0101110110101001    0101110110101010    0101110110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23975 - 23979

  --0101110110101100    0101110110101101    0101110110101110    0101110110101111    0101110110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23980 - 23984

  --0101110110110001    0101110110110010    0101110110110011    0101110110110100    0101110110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23985 - 23989

  --0101110110110110    0101110110110111    0101110110111000    0101110110111001    0101110110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23990 - 23994

  --0101110110111011    0101110110111100    0101110110111101    0101110110111110    0101110110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 23995 - 23999

  --0101110111000000    0101110111000001    0101110111000010    0101110111000011    0101110111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24000 - 24004

  --0101110111000101    0101110111000110    0101110111000111    0101110111001000    0101110111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24005 - 24009

  --0101110111001010    0101110111001011    0101110111001100    0101110111001101    0101110111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24010 - 24014

  --0101110111001111    0101110111010000    0101110111010001    0101110111010010    0101110111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24015 - 24019

  --0101110111010100    0101110111010101    0101110111010110    0101110111010111    0101110111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24020 - 24024

  --0101110111011001    0101110111011010    0101110111011011    0101110111011100    0101110111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24025 - 24029

  --0101110111011110    0101110111011111    0101110111100000    0101110111100001    0101110111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24030 - 24034

  --0101110111100011    0101110111100100    0101110111100101    0101110111100110    0101110111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24035 - 24039

  --0101110111101000    0101110111101001    0101110111101010    0101110111101011    0101110111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24040 - 24044

  --0101110111101101    0101110111101110    0101110111101111    0101110111110000    0101110111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24045 - 24049

  --0101110111110010    0101110111110011    0101110111110100    0101110111110101    0101110111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24050 - 24054

  --0101110111110111    0101110111111000    0101110111111001    0101110111111010    0101110111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24055 - 24059

  --0101110111111100    0101110111111101    0101110111111110    0101110111111111    0101111000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24060 - 24064

  --0101111000000001    0101111000000010    0101111000000011    0101111000000100    0101111000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24065 - 24069

  --0101111000000110    0101111000000111    0101111000001000    0101111000001001    0101111000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24070 - 24074

  --0101111000001011    0101111000001100    0101111000001101    0101111000001110    0101111000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24075 - 24079

  --0101111000010000    0101111000010001    0101111000010010    0101111000010011    0101111000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24080 - 24084

  --0101111000010101    0101111000010110    0101111000010111    0101111000011000    0101111000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24085 - 24089

  --0101111000011010    0101111000011011    0101111000011100    0101111000011101    0101111000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24090 - 24094

  --0101111000011111    0101111000100000    0101111000100001    0101111000100010    0101111000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24095 - 24099

  --0101111000100100    0101111000100101    0101111000100110    0101111000100111    0101111000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24100 - 24104

  --0101111000101001    0101111000101010    0101111000101011    0101111000101100    0101111000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24105 - 24109

  --0101111000101110    0101111000101111    0101111000110000    0101111000110001    0101111000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24110 - 24114

  --0101111000110011    0101111000110100    0101111000110101    0101111000110110    0101111000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24115 - 24119

  --0101111000111000    0101111000111001    0101111000111010    0101111000111011    0101111000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24120 - 24124

  --0101111000111101    0101111000111110    0101111000111111    0101111001000000    0101111001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24125 - 24129

  --0101111001000010    0101111001000011    0101111001000100    0101111001000101    0101111001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24130 - 24134

  --0101111001000111    0101111001001000    0101111001001001    0101111001001010    0101111001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24135 - 24139

  --0101111001001100    0101111001001101    0101111001001110    0101111001001111    0101111001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24140 - 24144

  --0101111001010001    0101111001010010    0101111001010011    0101111001010100    0101111001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24145 - 24149

  --0101111001010110    0101111001010111    0101111001011000    0101111001011001    0101111001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24150 - 24154

  --0101111001011011    0101111001011100    0101111001011101    0101111001011110    0101111001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24155 - 24159

  --0101111001100000    0101111001100001    0101111001100010    0101111001100011    0101111001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24160 - 24164

  --0101111001100101    0101111001100110    0101111001100111    0101111001101000    0101111001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24165 - 24169

  --0101111001101010    0101111001101011    0101111001101100    0101111001101101    0101111001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24170 - 24174

  --0101111001101111    0101111001110000    0101111001110001    0101111001110010    0101111001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24175 - 24179

  --0101111001110100    0101111001110101    0101111001110110    0101111001110111    0101111001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24180 - 24184

  --0101111001111001    0101111001111010    0101111001111011    0101111001111100    0101111001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24185 - 24189

  --0101111001111110    0101111001111111    0101111010000000    0101111010000001    0101111010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24190 - 24194

  --0101111010000011    0101111010000100    0101111010000101    0101111010000110    0101111010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24195 - 24199

  --0101111010001000    0101111010001001    0101111010001010    0101111010001011    0101111010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24200 - 24204

  --0101111010001101    0101111010001110    0101111010001111    0101111010010000    0101111010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24205 - 24209

  --0101111010010010    0101111010010011    0101111010010100    0101111010010101    0101111010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24210 - 24214

  --0101111010010111    0101111010011000    0101111010011001    0101111010011010    0101111010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24215 - 24219

  --0101111010011100    0101111010011101    0101111010011110    0101111010011111    0101111010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24220 - 24224

  --0101111010100001    0101111010100010    0101111010100011    0101111010100100    0101111010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24225 - 24229

  --0101111010100110    0101111010100111    0101111010101000    0101111010101001    0101111010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24230 - 24234

  --0101111010101011    0101111010101100    0101111010101101    0101111010101110    0101111010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24235 - 24239

  --0101111010110000    0101111010110001    0101111010110010    0101111010110011    0101111010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24240 - 24244

  --0101111010110101    0101111010110110    0101111010110111    0101111010111000    0101111010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24245 - 24249

  --0101111010111010    0101111010111011    0101111010111100    0101111010111101    0101111010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24250 - 24254

  --0101111010111111    0101111011000000    0101111011000001    0101111011000010    0101111011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24255 - 24259

  --0101111011000100    0101111011000101    0101111011000110    0101111011000111    0101111011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24260 - 24264

  --0101111011001001    0101111011001010    0101111011001011    0101111011001100    0101111011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24265 - 24269

  --0101111011001110    0101111011001111    0101111011010000    0101111011010001    0101111011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24270 - 24274

  --0101111011010011    0101111011010100    0101111011010101    0101111011010110    0101111011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24275 - 24279

  --0101111011011000    0101111011011001    0101111011011010    0101111011011011    0101111011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24280 - 24284

  --0101111011011101    0101111011011110    0101111011011111    0101111011100000    0101111011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24285 - 24289

  --0101111011100010    0101111011100011    0101111011100100    0101111011100101    0101111011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24290 - 24294

  --0101111011100111    0101111011101000    0101111011101001    0101111011101010    0101111011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24295 - 24299

  --0101111011101100    0101111011101101    0101111011101110    0101111011101111    0101111011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24300 - 24304

  --0101111011110001    0101111011110010    0101111011110011    0101111011110100    0101111011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24305 - 24309

  --0101111011110110    0101111011110111    0101111011111000    0101111011111001    0101111011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24310 - 24314

  --0101111011111011    0101111011111100    0101111011111101    0101111011111110    0101111011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24315 - 24319

  --0101111100000000    0101111100000001    0101111100000010    0101111100000011    0101111100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24320 - 24324

  --0101111100000101    0101111100000110    0101111100000111    0101111100001000    0101111100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24325 - 24329

  --0101111100001010    0101111100001011    0101111100001100    0101111100001101    0101111100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24330 - 24334

  --0101111100001111    0101111100010000    0101111100010001    0101111100010010    0101111100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24335 - 24339

  --0101111100010100    0101111100010101    0101111100010110    0101111100010111    0101111100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24340 - 24344

  --0101111100011001    0101111100011010    0101111100011011    0101111100011100    0101111100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24345 - 24349

  --0101111100011110    0101111100011111    0101111100100000    0101111100100001    0101111100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24350 - 24354

  --0101111100100011    0101111100100100    0101111100100101    0101111100100110    0101111100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24355 - 24359

  --0101111100101000    0101111100101001    0101111100101010    0101111100101011    0101111100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24360 - 24364

  --0101111100101101    0101111100101110    0101111100101111    0101111100110000    0101111100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24365 - 24369

  --0101111100110010    0101111100110011    0101111100110100    0101111100110101    0101111100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24370 - 24374

  --0101111100110111    0101111100111000    0101111100111001    0101111100111010    0101111100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24375 - 24379

  --0101111100111100    0101111100111101    0101111100111110    0101111100111111    0101111101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24380 - 24384

  --0101111101000001    0101111101000010    0101111101000011    0101111101000100    0101111101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24385 - 24389

  --0101111101000110    0101111101000111    0101111101001000    0101111101001001    0101111101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24390 - 24394

  --0101111101001011    0101111101001100    0101111101001101    0101111101001110    0101111101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24395 - 24399

  --0101111101010000    0101111101010001    0101111101010010    0101111101010011    0101111101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24400 - 24404

  --0101111101010101    0101111101010110    0101111101010111    0101111101011000    0101111101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24405 - 24409

  --0101111101011010    0101111101011011    0101111101011100    0101111101011101    0101111101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24410 - 24414

  --0101111101011111    0101111101100000    0101111101100001    0101111101100010    0101111101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24415 - 24419

  --0101111101100100    0101111101100101    0101111101100110    0101111101100111    0101111101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24420 - 24424

  --0101111101101001    0101111101101010    0101111101101011    0101111101101100    0101111101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24425 - 24429

  --0101111101101110    0101111101101111    0101111101110000    0101111101110001    0101111101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24430 - 24434

  --0101111101110011    0101111101110100    0101111101110101    0101111101110110    0101111101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24435 - 24439

  --0101111101111000    0101111101111001    0101111101111010    0101111101111011    0101111101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24440 - 24444

  --0101111101111101    0101111101111110    0101111101111111    0101111110000000    0101111110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24445 - 24449

  --0101111110000010    0101111110000011    0101111110000100    0101111110000101    0101111110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24450 - 24454

  --0101111110000111    0101111110001000    0101111110001001    0101111110001010    0101111110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24455 - 24459

  --0101111110001100    0101111110001101    0101111110001110    0101111110001111    0101111110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24460 - 24464

  --0101111110010001    0101111110010010    0101111110010011    0101111110010100    0101111110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24465 - 24469

  --0101111110010110    0101111110010111    0101111110011000    0101111110011001    0101111110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24470 - 24474

  --0101111110011011    0101111110011100    0101111110011101    0101111110011110    0101111110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24475 - 24479

  --0101111110100000    0101111110100001    0101111110100010    0101111110100011    0101111110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24480 - 24484

  --0101111110100101    0101111110100110    0101111110100111    0101111110101000    0101111110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24485 - 24489

  --0101111110101010    0101111110101011    0101111110101100    0101111110101101    0101111110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24490 - 24494

  --0101111110101111    0101111110110000    0101111110110001    0101111110110010    0101111110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24495 - 24499

  --0101111110110100    0101111110110101    0101111110110110    0101111110110111    0101111110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24500 - 24504

  --0101111110111001    0101111110111010    0101111110111011    0101111110111100    0101111110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24505 - 24509

  --0101111110111110    0101111110111111    0101111111000000    0101111111000001    0101111111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24510 - 24514

  --0101111111000011    0101111111000100    0101111111000101    0101111111000110    0101111111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24515 - 24519

  --0101111111001000    0101111111001001    0101111111001010    0101111111001011    0101111111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24520 - 24524

  --0101111111001101    0101111111001110    0101111111001111    0101111111010000    0101111111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24525 - 24529

  --0101111111010010    0101111111010011    0101111111010100    0101111111010101    0101111111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24530 - 24534

  --0101111111010111    0101111111011000    0101111111011001    0101111111011010    0101111111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24535 - 24539

  --0101111111011100    0101111111011101    0101111111011110    0101111111011111    0101111111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24540 - 24544

  --0101111111100001    0101111111100010    0101111111100011    0101111111100100    0101111111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24545 - 24549

  --0101111111100110    0101111111100111    0101111111101000    0101111111101001    0101111111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24550 - 24554

  --0101111111101011    0101111111101100    0101111111101101    0101111111101110    0101111111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24555 - 24559

  --0101111111110000    0101111111110001    0101111111110010    0101111111110011    0101111111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24560 - 24564

  --0101111111110101    0101111111110110    0101111111110111    0101111111111000    0101111111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24565 - 24569

  --0101111111111010    0101111111111011    0101111111111100    0101111111111101    0101111111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24570 - 24574

  --0101111111111111    0110000000000000    0110000000000001    0110000000000010    0110000000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24575 - 24579

  --0110000000000100    0110000000000101    0110000000000110    0110000000000111    0110000000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24580 - 24584

  --0110000000001001    0110000000001010    0110000000001011    0110000000001100    0110000000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24585 - 24589

  --0110000000001110    0110000000001111    0110000000010000    0110000000010001    0110000000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24590 - 24594

  --0110000000010011    0110000000010100    0110000000010101    0110000000010110    0110000000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24595 - 24599

  --0110000000011000    0110000000011001    0110000000011010    0110000000011011    0110000000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24600 - 24604

  --0110000000011101    0110000000011110    0110000000011111    0110000000100000    0110000000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24605 - 24609

  --0110000000100010    0110000000100011    0110000000100100    0110000000100101    0110000000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24610 - 24614

  --0110000000100111    0110000000101000    0110000000101001    0110000000101010    0110000000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24615 - 24619

  --0110000000101100    0110000000101101    0110000000101110    0110000000101111    0110000000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24620 - 24624

  --0110000000110001    0110000000110010    0110000000110011    0110000000110100    0110000000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24625 - 24629

  --0110000000110110    0110000000110111    0110000000111000    0110000000111001    0110000000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24630 - 24634

  --0110000000111011    0110000000111100    0110000000111101    0110000000111110    0110000000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24635 - 24639

  --0110000001000000    0110000001000001    0110000001000010    0110000001000011    0110000001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24640 - 24644

  --0110000001000101    0110000001000110    0110000001000111    0110000001001000    0110000001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24645 - 24649

  --0110000001001010    0110000001001011    0110000001001100    0110000001001101    0110000001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24650 - 24654

  --0110000001001111    0110000001010000    0110000001010001    0110000001010010    0110000001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24655 - 24659

  --0110000001010100    0110000001010101    0110000001010110    0110000001010111    0110000001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24660 - 24664

  --0110000001011001    0110000001011010    0110000001011011    0110000001011100    0110000001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24665 - 24669

  --0110000001011110    0110000001011111    0110000001100000    0110000001100001    0110000001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24670 - 24674

  --0110000001100011    0110000001100100    0110000001100101    0110000001100110    0110000001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24675 - 24679

  --0110000001101000    0110000001101001    0110000001101010    0110000001101011    0110000001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24680 - 24684

  --0110000001101101    0110000001101110    0110000001101111    0110000001110000    0110000001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24685 - 24689

  --0110000001110010    0110000001110011    0110000001110100    0110000001110101    0110000001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24690 - 24694

  --0110000001110111    0110000001111000    0110000001111001    0110000001111010    0110000001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24695 - 24699

  --0110000001111100    0110000001111101    0110000001111110    0110000001111111    0110000010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24700 - 24704

  --0110000010000001    0110000010000010    0110000010000011    0110000010000100    0110000010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24705 - 24709

  --0110000010000110    0110000010000111    0110000010001000    0110000010001001    0110000010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24710 - 24714

  --0110000010001011    0110000010001100    0110000010001101    0110000010001110    0110000010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24715 - 24719

  --0110000010010000    0110000010010001    0110000010010010    0110000010010011    0110000010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24720 - 24724

  --0110000010010101    0110000010010110    0110000010010111    0110000010011000    0110000010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24725 - 24729

  --0110000010011010    0110000010011011    0110000010011100    0110000010011101    0110000010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24730 - 24734

  --0110000010011111    0110000010100000    0110000010100001    0110000010100010    0110000010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24735 - 24739

  --0110000010100100    0110000010100101    0110000010100110    0110000010100111    0110000010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24740 - 24744

  --0110000010101001    0110000010101010    0110000010101011    0110000010101100    0110000010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24745 - 24749

  --0110000010101110    0110000010101111    0110000010110000    0110000010110001    0110000010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24750 - 24754

  --0110000010110011    0110000010110100    0110000010110101    0110000010110110    0110000010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24755 - 24759

  --0110000010111000    0110000010111001    0110000010111010    0110000010111011    0110000010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24760 - 24764

  --0110000010111101    0110000010111110    0110000010111111    0110000011000000    0110000011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24765 - 24769

  --0110000011000010    0110000011000011    0110000011000100    0110000011000101    0110000011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24770 - 24774

  --0110000011000111    0110000011001000    0110000011001001    0110000011001010    0110000011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24775 - 24779

  --0110000011001100    0110000011001101    0110000011001110    0110000011001111    0110000011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24780 - 24784

  --0110000011010001    0110000011010010    0110000011010011    0110000011010100    0110000011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24785 - 24789

  --0110000011010110    0110000011010111    0110000011011000    0110000011011001    0110000011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24790 - 24794

  --0110000011011011    0110000011011100    0110000011011101    0110000011011110    0110000011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24795 - 24799

  --0110000011100000    0110000011100001    0110000011100010    0110000011100011    0110000011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24800 - 24804

  --0110000011100101    0110000011100110    0110000011100111    0110000011101000    0110000011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24805 - 24809

  --0110000011101010    0110000011101011    0110000011101100    0110000011101101    0110000011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24810 - 24814

  --0110000011101111    0110000011110000    0110000011110001    0110000011110010    0110000011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24815 - 24819

  --0110000011110100    0110000011110101    0110000011110110    0110000011110111    0110000011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24820 - 24824

  --0110000011111001    0110000011111010    0110000011111011    0110000011111100    0110000011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24825 - 24829

  --0110000011111110    0110000011111111    0110000100000000    0110000100000001    0110000100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24830 - 24834

  --0110000100000011    0110000100000100    0110000100000101    0110000100000110    0110000100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24835 - 24839

  --0110000100001000    0110000100001001    0110000100001010    0110000100001011    0110000100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24840 - 24844

  --0110000100001101    0110000100001110    0110000100001111    0110000100010000    0110000100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24845 - 24849

  --0110000100010010    0110000100010011    0110000100010100    0110000100010101    0110000100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24850 - 24854

  --0110000100010111    0110000100011000    0110000100011001    0110000100011010    0110000100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24855 - 24859

  --0110000100011100    0110000100011101    0110000100011110    0110000100011111    0110000100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24860 - 24864

  --0110000100100001    0110000100100010    0110000100100011    0110000100100100    0110000100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24865 - 24869

  --0110000100100110    0110000100100111    0110000100101000    0110000100101001    0110000100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24870 - 24874

  --0110000100101011    0110000100101100    0110000100101101    0110000100101110    0110000100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24875 - 24879

  --0110000100110000    0110000100110001    0110000100110010    0110000100110011    0110000100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24880 - 24884

  --0110000100110101    0110000100110110    0110000100110111    0110000100111000    0110000100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24885 - 24889

  --0110000100111010    0110000100111011    0110000100111100    0110000100111101    0110000100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24890 - 24894

  --0110000100111111    0110000101000000    0110000101000001    0110000101000010    0110000101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24895 - 24899

  --0110000101000100    0110000101000101    0110000101000110    0110000101000111    0110000101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24900 - 24904

  --0110000101001001    0110000101001010    0110000101001011    0110000101001100    0110000101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24905 - 24909

  --0110000101001110    0110000101001111    0110000101010000    0110000101010001    0110000101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24910 - 24914

  --0110000101010011    0110000101010100    0110000101010101    0110000101010110    0110000101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24915 - 24919

  --0110000101011000    0110000101011001    0110000101011010    0110000101011011    0110000101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24920 - 24924

  --0110000101011101    0110000101011110    0110000101011111    0110000101100000    0110000101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24925 - 24929

  --0110000101100010    0110000101100011    0110000101100100    0110000101100101    0110000101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24930 - 24934

  --0110000101100111    0110000101101000    0110000101101001    0110000101101010    0110000101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24935 - 24939

  --0110000101101100    0110000101101101    0110000101101110    0110000101101111    0110000101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24940 - 24944

  --0110000101110001    0110000101110010    0110000101110011    0110000101110100    0110000101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24945 - 24949

  --0110000101110110    0110000101110111    0110000101111000    0110000101111001    0110000101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24950 - 24954

  --0110000101111011    0110000101111100    0110000101111101    0110000101111110    0110000101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24955 - 24959

  --0110000110000000    0110000110000001    0110000110000010    0110000110000011    0110000110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24960 - 24964

  --0110000110000101    0110000110000110    0110000110000111    0110000110001000    0110000110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24965 - 24969

  --0110000110001010    0110000110001011    0110000110001100    0110000110001101    0110000110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24970 - 24974

  --0110000110001111    0110000110010000    0110000110010001    0110000110010010    0110000110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24975 - 24979

  --0110000110010100    0110000110010101    0110000110010110    0110000110010111    0110000110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24980 - 24984

  --0110000110011001    0110000110011010    0110000110011011    0110000110011100    0110000110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24985 - 24989

  --0110000110011110    0110000110011111    0110000110100000    0110000110100001    0110000110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24990 - 24994

  --0110000110100011    0110000110100100    0110000110100101    0110000110100110    0110000110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 24995 - 24999

  --0110000110101000    0110000110101001    0110000110101010    0110000110101011    0110000110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25000 - 25004

  --0110000110101101    0110000110101110    0110000110101111    0110000110110000    0110000110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25005 - 25009

  --0110000110110010    0110000110110011    0110000110110100    0110000110110101    0110000110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25010 - 25014

  --0110000110110111    0110000110111000    0110000110111001    0110000110111010    0110000110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25015 - 25019

  --0110000110111100    0110000110111101    0110000110111110    0110000110111111    0110000111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25020 - 25024

  --0110000111000001    0110000111000010    0110000111000011    0110000111000100    0110000111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25025 - 25029

  --0110000111000110    0110000111000111    0110000111001000    0110000111001001    0110000111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25030 - 25034

  --0110000111001011    0110000111001100    0110000111001101    0110000111001110    0110000111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25035 - 25039

  --0110000111010000    0110000111010001    0110000111010010    0110000111010011    0110000111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25040 - 25044

  --0110000111010101    0110000111010110    0110000111010111    0110000111011000    0110000111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25045 - 25049

  --0110000111011010    0110000111011011    0110000111011100    0110000111011101    0110000111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25050 - 25054

  --0110000111011111    0110000111100000    0110000111100001    0110000111100010    0110000111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25055 - 25059

  --0110000111100100    0110000111100101    0110000111100110    0110000111100111    0110000111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25060 - 25064

  --0110000111101001    0110000111101010    0110000111101011    0110000111101100    0110000111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25065 - 25069

  --0110000111101110    0110000111101111    0110000111110000    0110000111110001    0110000111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25070 - 25074

  --0110000111110011    0110000111110100    0110000111110101    0110000111110110    0110000111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25075 - 25079

  --0110000111111000    0110000111111001    0110000111111010    0110000111111011    0110000111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25080 - 25084

  --0110000111111101    0110000111111110    0110000111111111    0110001000000000    0110001000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25085 - 25089

  --0110001000000010    0110001000000011    0110001000000100    0110001000000101    0110001000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25090 - 25094

  --0110001000000111    0110001000001000    0110001000001001    0110001000001010    0110001000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25095 - 25099

  --0110001000001100    0110001000001101    0110001000001110    0110001000001111    0110001000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25100 - 25104

  --0110001000010001    0110001000010010    0110001000010011    0110001000010100    0110001000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25105 - 25109

  --0110001000010110    0110001000010111    0110001000011000    0110001000011001    0110001000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25110 - 25114

  --0110001000011011    0110001000011100    0110001000011101    0110001000011110    0110001000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25115 - 25119

  --0110001000100000    0110001000100001    0110001000100010    0110001000100011    0110001000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25120 - 25124

  --0110001000100101    0110001000100110    0110001000100111    0110001000101000    0110001000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25125 - 25129

  --0110001000101010    0110001000101011    0110001000101100    0110001000101101    0110001000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25130 - 25134

  --0110001000101111    0110001000110000    0110001000110001    0110001000110010    0110001000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25135 - 25139

  --0110001000110100    0110001000110101    0110001000110110    0110001000110111    0110001000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25140 - 25144

  --0110001000111001    0110001000111010    0110001000111011    0110001000111100    0110001000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25145 - 25149

  --0110001000111110    0110001000111111    0110001001000000    0110001001000001    0110001001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25150 - 25154

  --0110001001000011    0110001001000100    0110001001000101    0110001001000110    0110001001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25155 - 25159

  --0110001001001000    0110001001001001    0110001001001010    0110001001001011    0110001001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25160 - 25164

  --0110001001001101    0110001001001110    0110001001001111    0110001001010000    0110001001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25165 - 25169

  --0110001001010010    0110001001010011    0110001001010100    0110001001010101    0110001001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25170 - 25174

  --0110001001010111    0110001001011000    0110001001011001    0110001001011010    0110001001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25175 - 25179

  --0110001001011100    0110001001011101    0110001001011110    0110001001011111    0110001001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25180 - 25184

  --0110001001100001    0110001001100010    0110001001100011    0110001001100100    0110001001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25185 - 25189

  --0110001001100110    0110001001100111    0110001001101000    0110001001101001    0110001001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25190 - 25194

  --0110001001101011    0110001001101100    0110001001101101    0110001001101110    0110001001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25195 - 25199

  --0110001001110000    0110001001110001    0110001001110010    0110001001110011    0110001001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25200 - 25204

  --0110001001110101    0110001001110110    0110001001110111    0110001001111000    0110001001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25205 - 25209

  --0110001001111010    0110001001111011    0110001001111100    0110001001111101    0110001001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25210 - 25214

  --0110001001111111    0110001010000000    0110001010000001    0110001010000010    0110001010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25215 - 25219

  --0110001010000100    0110001010000101    0110001010000110    0110001010000111    0110001010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25220 - 25224

  --0110001010001001    0110001010001010    0110001010001011    0110001010001100    0110001010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25225 - 25229

  --0110001010001110    0110001010001111    0110001010010000    0110001010010001    0110001010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25230 - 25234

  --0110001010010011    0110001010010100    0110001010010101    0110001010010110    0110001010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25235 - 25239

  --0110001010011000    0110001010011001    0110001010011010    0110001010011011    0110001010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25240 - 25244

  --0110001010011101    0110001010011110    0110001010011111    0110001010100000    0110001010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25245 - 25249

  --0110001010100010    0110001010100011    0110001010100100    0110001010100101    0110001010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25250 - 25254

  --0110001010100111    0110001010101000    0110001010101001    0110001010101010    0110001010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25255 - 25259

  --0110001010101100    0110001010101101    0110001010101110    0110001010101111    0110001010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25260 - 25264

  --0110001010110001    0110001010110010    0110001010110011    0110001010110100    0110001010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25265 - 25269

  --0110001010110110    0110001010110111    0110001010111000    0110001010111001    0110001010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25270 - 25274

  --0110001010111011    0110001010111100    0110001010111101    0110001010111110    0110001010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25275 - 25279

  --0110001011000000    0110001011000001    0110001011000010    0110001011000011    0110001011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25280 - 25284

  --0110001011000101    0110001011000110    0110001011000111    0110001011001000    0110001011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25285 - 25289

  --0110001011001010    0110001011001011    0110001011001100    0110001011001101    0110001011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25290 - 25294

  --0110001011001111    0110001011010000    0110001011010001    0110001011010010    0110001011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25295 - 25299

  --0110001011010100    0110001011010101    0110001011010110    0110001011010111    0110001011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25300 - 25304

  --0110001011011001    0110001011011010    0110001011011011    0110001011011100    0110001011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25305 - 25309

  --0110001011011110    0110001011011111    0110001011100000    0110001011100001    0110001011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25310 - 25314

  --0110001011100011    0110001011100100    0110001011100101    0110001011100110    0110001011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25315 - 25319

  --0110001011101000    0110001011101001    0110001011101010    0110001011101011    0110001011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25320 - 25324

  --0110001011101101    0110001011101110    0110001011101111    0110001011110000    0110001011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25325 - 25329

  --0110001011110010    0110001011110011    0110001011110100    0110001011110101    0110001011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25330 - 25334

  --0110001011110111    0110001011111000    0110001011111001    0110001011111010    0110001011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25335 - 25339

  --0110001011111100    0110001011111101    0110001011111110    0110001011111111    0110001100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25340 - 25344

  --0110001100000001    0110001100000010    0110001100000011    0110001100000100    0110001100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25345 - 25349

  --0110001100000110    0110001100000111    0110001100001000    0110001100001001    0110001100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25350 - 25354

  --0110001100001011    0110001100001100    0110001100001101    0110001100001110    0110001100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25355 - 25359

  --0110001100010000    0110001100010001    0110001100010010    0110001100010011    0110001100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25360 - 25364

  --0110001100010101    0110001100010110    0110001100010111    0110001100011000    0110001100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25365 - 25369

  --0110001100011010    0110001100011011    0110001100011100    0110001100011101    0110001100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25370 - 25374

  --0110001100011111    0110001100100000    0110001100100001    0110001100100010    0110001100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25375 - 25379

  --0110001100100100    0110001100100101    0110001100100110    0110001100100111    0110001100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25380 - 25384

  --0110001100101001    0110001100101010    0110001100101011    0110001100101100    0110001100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25385 - 25389

  --0110001100101110    0110001100101111    0110001100110000    0110001100110001    0110001100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25390 - 25394

  --0110001100110011    0110001100110100    0110001100110101    0110001100110110    0110001100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25395 - 25399

  --0110001100111000    0110001100111001    0110001100111010    0110001100111011    0110001100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25400 - 25404

  --0110001100111101    0110001100111110    0110001100111111    0110001101000000    0110001101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25405 - 25409

  --0110001101000010    0110001101000011    0110001101000100    0110001101000101    0110001101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25410 - 25414

  --0110001101000111    0110001101001000    0110001101001001    0110001101001010    0110001101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25415 - 25419

  --0110001101001100    0110001101001101    0110001101001110    0110001101001111    0110001101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25420 - 25424

  --0110001101010001    0110001101010010    0110001101010011    0110001101010100    0110001101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25425 - 25429

  --0110001101010110    0110001101010111    0110001101011000    0110001101011001    0110001101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25430 - 25434

  --0110001101011011    0110001101011100    0110001101011101    0110001101011110    0110001101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25435 - 25439

  --0110001101100000    0110001101100001    0110001101100010    0110001101100011    0110001101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25440 - 25444

  --0110001101100101    0110001101100110    0110001101100111    0110001101101000    0110001101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25445 - 25449

  --0110001101101010    0110001101101011    0110001101101100    0110001101101101    0110001101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25450 - 25454

  --0110001101101111    0110001101110000    0110001101110001    0110001101110010    0110001101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25455 - 25459

  --0110001101110100    0110001101110101    0110001101110110    0110001101110111    0110001101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25460 - 25464

  --0110001101111001    0110001101111010    0110001101111011    0110001101111100    0110001101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25465 - 25469

  --0110001101111110    0110001101111111    0110001110000000    0110001110000001    0110001110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25470 - 25474

  --0110001110000011    0110001110000100    0110001110000101    0110001110000110    0110001110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25475 - 25479

  --0110001110001000    0110001110001001    0110001110001010    0110001110001011    0110001110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25480 - 25484

  --0110001110001101    0110001110001110    0110001110001111    0110001110010000    0110001110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25485 - 25489

  --0110001110010010    0110001110010011    0110001110010100    0110001110010101    0110001110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25490 - 25494

  --0110001110010111    0110001110011000    0110001110011001    0110001110011010    0110001110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25495 - 25499

  --0110001110011100    0110001110011101    0110001110011110    0110001110011111    0110001110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25500 - 25504

  --0110001110100001    0110001110100010    0110001110100011    0110001110100100    0110001110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25505 - 25509

  --0110001110100110    0110001110100111    0110001110101000    0110001110101001    0110001110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25510 - 25514

  --0110001110101011    0110001110101100    0110001110101101    0110001110101110    0110001110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25515 - 25519

  --0110001110110000    0110001110110001    0110001110110010    0110001110110011    0110001110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25520 - 25524

  --0110001110110101    0110001110110110    0110001110110111    0110001110111000    0110001110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25525 - 25529

  --0110001110111010    0110001110111011    0110001110111100    0110001110111101    0110001110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25530 - 25534

  --0110001110111111    0110001111000000    0110001111000001    0110001111000010    0110001111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25535 - 25539

  --0110001111000100    0110001111000101    0110001111000110    0110001111000111    0110001111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25540 - 25544

  --0110001111001001    0110001111001010    0110001111001011    0110001111001100    0110001111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25545 - 25549

  --0110001111001110    0110001111001111    0110001111010000    0110001111010001    0110001111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25550 - 25554

  --0110001111010011    0110001111010100    0110001111010101    0110001111010110    0110001111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25555 - 25559

  --0110001111011000    0110001111011001    0110001111011010    0110001111011011    0110001111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25560 - 25564

  --0110001111011101    0110001111011110    0110001111011111    0110001111100000    0110001111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25565 - 25569

  --0110001111100010    0110001111100011    0110001111100100    0110001111100101    0110001111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25570 - 25574

  --0110001111100111    0110001111101000    0110001111101001    0110001111101010    0110001111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25575 - 25579

  --0110001111101100    0110001111101101    0110001111101110    0110001111101111    0110001111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25580 - 25584

  --0110001111110001    0110001111110010    0110001111110011    0110001111110100    0110001111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25585 - 25589

  --0110001111110110    0110001111110111    0110001111111000    0110001111111001    0110001111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25590 - 25594

  --0110001111111011    0110001111111100    0110001111111101    0110001111111110    0110001111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25595 - 25599

  --0110010000000000    0110010000000001    0110010000000010    0110010000000011    0110010000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25600 - 25604

  --0110010000000101    0110010000000110    0110010000000111    0110010000001000    0110010000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25605 - 25609

  --0110010000001010    0110010000001011    0110010000001100    0110010000001101    0110010000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25610 - 25614

  --0110010000001111    0110010000010000    0110010000010001    0110010000010010    0110010000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25615 - 25619

  --0110010000010100    0110010000010101    0110010000010110    0110010000010111    0110010000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25620 - 25624

  --0110010000011001    0110010000011010    0110010000011011    0110010000011100    0110010000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25625 - 25629

  --0110010000011110    0110010000011111    0110010000100000    0110010000100001    0110010000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25630 - 25634

  --0110010000100011    0110010000100100    0110010000100101    0110010000100110    0110010000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25635 - 25639

  --0110010000101000    0110010000101001    0110010000101010    0110010000101011    0110010000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25640 - 25644

  --0110010000101101    0110010000101110    0110010000101111    0110010000110000    0110010000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25645 - 25649

  --0110010000110010    0110010000110011    0110010000110100    0110010000110101    0110010000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25650 - 25654

  --0110010000110111    0110010000111000    0110010000111001    0110010000111010    0110010000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25655 - 25659

  --0110010000111100    0110010000111101    0110010000111110    0110010000111111    0110010001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25660 - 25664

  --0110010001000001    0110010001000010    0110010001000011    0110010001000100    0110010001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25665 - 25669

  --0110010001000110    0110010001000111    0110010001001000    0110010001001001    0110010001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25670 - 25674

  --0110010001001011    0110010001001100    0110010001001101    0110010001001110    0110010001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25675 - 25679

  --0110010001010000    0110010001010001    0110010001010010    0110010001010011    0110010001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25680 - 25684

  --0110010001010101    0110010001010110    0110010001010111    0110010001011000    0110010001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25685 - 25689

  --0110010001011010    0110010001011011    0110010001011100    0110010001011101    0110010001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25690 - 25694

  --0110010001011111    0110010001100000    0110010001100001    0110010001100010    0110010001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25695 - 25699

  --0110010001100100    0110010001100101    0110010001100110    0110010001100111    0110010001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25700 - 25704

  --0110010001101001    0110010001101010    0110010001101011    0110010001101100    0110010001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25705 - 25709

  --0110010001101110    0110010001101111    0110010001110000    0110010001110001    0110010001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25710 - 25714

  --0110010001110011    0110010001110100    0110010001110101    0110010001110110    0110010001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25715 - 25719

  --0110010001111000    0110010001111001    0110010001111010    0110010001111011    0110010001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25720 - 25724

  --0110010001111101    0110010001111110    0110010001111111    0110010010000000    0110010010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25725 - 25729

  --0110010010000010    0110010010000011    0110010010000100    0110010010000101    0110010010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25730 - 25734

  --0110010010000111    0110010010001000    0110010010001001    0110010010001010    0110010010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25735 - 25739

  --0110010010001100    0110010010001101    0110010010001110    0110010010001111    0110010010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25740 - 25744

  --0110010010010001    0110010010010010    0110010010010011    0110010010010100    0110010010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25745 - 25749

  --0110010010010110    0110010010010111    0110010010011000    0110010010011001    0110010010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25750 - 25754

  --0110010010011011    0110010010011100    0110010010011101    0110010010011110    0110010010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25755 - 25759

  --0110010010100000    0110010010100001    0110010010100010    0110010010100011    0110010010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25760 - 25764

  --0110010010100101    0110010010100110    0110010010100111    0110010010101000    0110010010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25765 - 25769

  --0110010010101010    0110010010101011    0110010010101100    0110010010101101    0110010010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25770 - 25774

  --0110010010101111    0110010010110000    0110010010110001    0110010010110010    0110010010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25775 - 25779

  --0110010010110100    0110010010110101    0110010010110110    0110010010110111    0110010010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25780 - 25784

  --0110010010111001    0110010010111010    0110010010111011    0110010010111100    0110010010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25785 - 25789

  --0110010010111110    0110010010111111    0110010011000000    0110010011000001    0110010011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25790 - 25794

  --0110010011000011    0110010011000100    0110010011000101    0110010011000110    0110010011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25795 - 25799

  --0110010011001000    0110010011001001    0110010011001010    0110010011001011    0110010011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25800 - 25804

  --0110010011001101    0110010011001110    0110010011001111    0110010011010000    0110010011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25805 - 25809

  --0110010011010010    0110010011010011    0110010011010100    0110010011010101    0110010011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25810 - 25814

  --0110010011010111    0110010011011000    0110010011011001    0110010011011010    0110010011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25815 - 25819

  --0110010011011100    0110010011011101    0110010011011110    0110010011011111    0110010011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25820 - 25824

  --0110010011100001    0110010011100010    0110010011100011    0110010011100100    0110010011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25825 - 25829

  --0110010011100110    0110010011100111    0110010011101000    0110010011101001    0110010011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25830 - 25834

  --0110010011101011    0110010011101100    0110010011101101    0110010011101110    0110010011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25835 - 25839

  --0110010011110000    0110010011110001    0110010011110010    0110010011110011    0110010011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25840 - 25844

  --0110010011110101    0110010011110110    0110010011110111    0110010011111000    0110010011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25845 - 25849

  --0110010011111010    0110010011111011    0110010011111100    0110010011111101    0110010011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25850 - 25854

  --0110010011111111    0110010100000000    0110010100000001    0110010100000010    0110010100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25855 - 25859

  --0110010100000100    0110010100000101    0110010100000110    0110010100000111    0110010100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25860 - 25864

  --0110010100001001    0110010100001010    0110010100001011    0110010100001100    0110010100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25865 - 25869

  --0110010100001110    0110010100001111    0110010100010000    0110010100010001    0110010100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25870 - 25874

  --0110010100010011    0110010100010100    0110010100010101    0110010100010110    0110010100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25875 - 25879

  --0110010100011000    0110010100011001    0110010100011010    0110010100011011    0110010100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25880 - 25884

  --0110010100011101    0110010100011110    0110010100011111    0110010100100000    0110010100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25885 - 25889

  --0110010100100010    0110010100100011    0110010100100100    0110010100100101    0110010100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25890 - 25894

  --0110010100100111    0110010100101000    0110010100101001    0110010100101010    0110010100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25895 - 25899

  --0110010100101100    0110010100101101    0110010100101110    0110010100101111    0110010100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25900 - 25904

  --0110010100110001    0110010100110010    0110010100110011    0110010100110100    0110010100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25905 - 25909

  --0110010100110110    0110010100110111    0110010100111000    0110010100111001    0110010100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25910 - 25914

  --0110010100111011    0110010100111100    0110010100111101    0110010100111110    0110010100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25915 - 25919

  --0110010101000000    0110010101000001    0110010101000010    0110010101000011    0110010101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25920 - 25924

  --0110010101000101    0110010101000110    0110010101000111    0110010101001000    0110010101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25925 - 25929

  --0110010101001010    0110010101001011    0110010101001100    0110010101001101    0110010101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25930 - 25934

  --0110010101001111    0110010101010000    0110010101010001    0110010101010010    0110010101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25935 - 25939

  --0110010101010100    0110010101010101    0110010101010110    0110010101010111    0110010101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25940 - 25944

  --0110010101011001    0110010101011010    0110010101011011    0110010101011100    0110010101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25945 - 25949

  --0110010101011110    0110010101011111    0110010101100000    0110010101100001    0110010101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25950 - 25954

  --0110010101100011    0110010101100100    0110010101100101    0110010101100110    0110010101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25955 - 25959

  --0110010101101000    0110010101101001    0110010101101010    0110010101101011    0110010101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25960 - 25964

  --0110010101101101    0110010101101110    0110010101101111    0110010101110000    0110010101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25965 - 25969

  --0110010101110010    0110010101110011    0110010101110100    0110010101110101    0110010101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25970 - 25974

  --0110010101110111    0110010101111000    0110010101111001    0110010101111010    0110010101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25975 - 25979

  --0110010101111100    0110010101111101    0110010101111110    0110010101111111    0110010110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25980 - 25984

  --0110010110000001    0110010110000010    0110010110000011    0110010110000100    0110010110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25985 - 25989

  --0110010110000110    0110010110000111    0110010110001000    0110010110001001    0110010110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25990 - 25994

  --0110010110001011    0110010110001100    0110010110001101    0110010110001110    0110010110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 25995 - 25999

  --0110010110010000    0110010110010001    0110010110010010    0110010110010011    0110010110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26000 - 26004

  --0110010110010101    0110010110010110    0110010110010111    0110010110011000    0110010110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26005 - 26009

  --0110010110011010    0110010110011011    0110010110011100    0110010110011101    0110010110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26010 - 26014

  --0110010110011111    0110010110100000    0110010110100001    0110010110100010    0110010110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26015 - 26019

  --0110010110100100    0110010110100101    0110010110100110    0110010110100111    0110010110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26020 - 26024

  --0110010110101001    0110010110101010    0110010110101011    0110010110101100    0110010110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26025 - 26029

  --0110010110101110    0110010110101111    0110010110110000    0110010110110001    0110010110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26030 - 26034

  --0110010110110011    0110010110110100    0110010110110101    0110010110110110    0110010110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26035 - 26039

  --0110010110111000    0110010110111001    0110010110111010    0110010110111011    0110010110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26040 - 26044

  --0110010110111101    0110010110111110    0110010110111111    0110010111000000    0110010111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26045 - 26049

  --0110010111000010    0110010111000011    0110010111000100    0110010111000101    0110010111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26050 - 26054

  --0110010111000111    0110010111001000    0110010111001001    0110010111001010    0110010111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26055 - 26059

  --0110010111001100    0110010111001101    0110010111001110    0110010111001111    0110010111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26060 - 26064

  --0110010111010001    0110010111010010    0110010111010011    0110010111010100    0110010111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26065 - 26069

  --0110010111010110    0110010111010111    0110010111011000    0110010111011001    0110010111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26070 - 26074

  --0110010111011011    0110010111011100    0110010111011101    0110010111011110    0110010111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26075 - 26079

  --0110010111100000    0110010111100001    0110010111100010    0110010111100011    0110010111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26080 - 26084

  --0110010111100101    0110010111100110    0110010111100111    0110010111101000    0110010111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26085 - 26089

  --0110010111101010    0110010111101011    0110010111101100    0110010111101101    0110010111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26090 - 26094

  --0110010111101111    0110010111110000    0110010111110001    0110010111110010    0110010111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26095 - 26099

  --0110010111110100    0110010111110101    0110010111110110    0110010111110111    0110010111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26100 - 26104

  --0110010111111001    0110010111111010    0110010111111011    0110010111111100    0110010111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26105 - 26109

  --0110010111111110    0110010111111111    0110011000000000    0110011000000001    0110011000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26110 - 26114

  --0110011000000011    0110011000000100    0110011000000101    0110011000000110    0110011000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26115 - 26119

  --0110011000001000    0110011000001001    0110011000001010    0110011000001011    0110011000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26120 - 26124

  --0110011000001101    0110011000001110    0110011000001111    0110011000010000    0110011000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26125 - 26129

  --0110011000010010    0110011000010011    0110011000010100    0110011000010101    0110011000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26130 - 26134

  --0110011000010111    0110011000011000    0110011000011001    0110011000011010    0110011000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26135 - 26139

  --0110011000011100    0110011000011101    0110011000011110    0110011000011111    0110011000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26140 - 26144

  --0110011000100001    0110011000100010    0110011000100011    0110011000100100    0110011000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26145 - 26149

  --0110011000100110    0110011000100111    0110011000101000    0110011000101001    0110011000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26150 - 26154

  --0110011000101011    0110011000101100    0110011000101101    0110011000101110    0110011000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26155 - 26159

  --0110011000110000    0110011000110001    0110011000110010    0110011000110011    0110011000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26160 - 26164

  --0110011000110101    0110011000110110    0110011000110111    0110011000111000    0110011000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26165 - 26169

  --0110011000111010    0110011000111011    0110011000111100    0110011000111101    0110011000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26170 - 26174

  --0110011000111111    0110011001000000    0110011001000001    0110011001000010    0110011001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26175 - 26179

  --0110011001000100    0110011001000101    0110011001000110    0110011001000111    0110011001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26180 - 26184

  --0110011001001001    0110011001001010    0110011001001011    0110011001001100    0110011001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26185 - 26189

  --0110011001001110    0110011001001111    0110011001010000    0110011001010001    0110011001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26190 - 26194

  --0110011001010011    0110011001010100    0110011001010101    0110011001010110    0110011001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26195 - 26199

  --0110011001011000    0110011001011001    0110011001011010    0110011001011011    0110011001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26200 - 26204

  --0110011001011101    0110011001011110    0110011001011111    0110011001100000    0110011001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26205 - 26209

  --0110011001100010    0110011001100011    0110011001100100    0110011001100101    0110011001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26210 - 26214

  --0110011001100111    0110011001101000    0110011001101001    0110011001101010    0110011001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26215 - 26219

  --0110011001101100    0110011001101101    0110011001101110    0110011001101111    0110011001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26220 - 26224

  --0110011001110001    0110011001110010    0110011001110011    0110011001110100    0110011001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26225 - 26229

  --0110011001110110    0110011001110111    0110011001111000    0110011001111001    0110011001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26230 - 26234

  --0110011001111011    0110011001111100    0110011001111101    0110011001111110    0110011001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26235 - 26239

  --0110011010000000    0110011010000001    0110011010000010    0110011010000011    0110011010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26240 - 26244

  --0110011010000101    0110011010000110    0110011010000111    0110011010001000    0110011010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26245 - 26249

  --0110011010001010    0110011010001011    0110011010001100    0110011010001101    0110011010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26250 - 26254

  --0110011010001111    0110011010010000    0110011010010001    0110011010010010    0110011010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26255 - 26259

  --0110011010010100    0110011010010101    0110011010010110    0110011010010111    0110011010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26260 - 26264

  --0110011010011001    0110011010011010    0110011010011011    0110011010011100    0110011010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26265 - 26269

  --0110011010011110    0110011010011111    0110011010100000    0110011010100001    0110011010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26270 - 26274

  --0110011010100011    0110011010100100    0110011010100101    0110011010100110    0110011010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26275 - 26279

  --0110011010101000    0110011010101001    0110011010101010    0110011010101011    0110011010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26280 - 26284

  --0110011010101101    0110011010101110    0110011010101111    0110011010110000    0110011010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26285 - 26289

  --0110011010110010    0110011010110011    0110011010110100    0110011010110101    0110011010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26290 - 26294

  --0110011010110111    0110011010111000    0110011010111001    0110011010111010    0110011010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26295 - 26299

  --0110011010111100    0110011010111101    0110011010111110    0110011010111111    0110011011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26300 - 26304

  --0110011011000001    0110011011000010    0110011011000011    0110011011000100    0110011011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26305 - 26309

  --0110011011000110    0110011011000111    0110011011001000    0110011011001001    0110011011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26310 - 26314

  --0110011011001011    0110011011001100    0110011011001101    0110011011001110    0110011011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26315 - 26319

  --0110011011010000    0110011011010001    0110011011010010    0110011011010011    0110011011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26320 - 26324

  --0110011011010101    0110011011010110    0110011011010111    0110011011011000    0110011011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26325 - 26329

  --0110011011011010    0110011011011011    0110011011011100    0110011011011101    0110011011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26330 - 26334

  --0110011011011111    0110011011100000    0110011011100001    0110011011100010    0110011011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26335 - 26339

  --0110011011100100    0110011011100101    0110011011100110    0110011011100111    0110011011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26340 - 26344

  --0110011011101001    0110011011101010    0110011011101011    0110011011101100    0110011011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26345 - 26349

  --0110011011101110    0110011011101111    0110011011110000    0110011011110001    0110011011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26350 - 26354

  --0110011011110011    0110011011110100    0110011011110101    0110011011110110    0110011011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26355 - 26359

  --0110011011111000    0110011011111001    0110011011111010    0110011011111011    0110011011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26360 - 26364

  --0110011011111101    0110011011111110    0110011011111111    0110011100000000    0110011100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26365 - 26369

  --0110011100000010    0110011100000011    0110011100000100    0110011100000101    0110011100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26370 - 26374

  --0110011100000111    0110011100001000    0110011100001001    0110011100001010    0110011100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26375 - 26379

  --0110011100001100    0110011100001101    0110011100001110    0110011100001111    0110011100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26380 - 26384

  --0110011100010001    0110011100010010    0110011100010011    0110011100010100    0110011100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26385 - 26389

  --0110011100010110    0110011100010111    0110011100011000    0110011100011001    0110011100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26390 - 26394

  --0110011100011011    0110011100011100    0110011100011101    0110011100011110    0110011100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26395 - 26399

  --0110011100100000    0110011100100001    0110011100100010    0110011100100011    0110011100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26400 - 26404

  --0110011100100101    0110011100100110    0110011100100111    0110011100101000    0110011100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26405 - 26409

  --0110011100101010    0110011100101011    0110011100101100    0110011100101101    0110011100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26410 - 26414

  --0110011100101111    0110011100110000    0110011100110001    0110011100110010    0110011100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26415 - 26419

  --0110011100110100    0110011100110101    0110011100110110    0110011100110111    0110011100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26420 - 26424

  --0110011100111001    0110011100111010    0110011100111011    0110011100111100    0110011100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26425 - 26429

  --0110011100111110    0110011100111111    0110011101000000    0110011101000001    0110011101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26430 - 26434

  --0110011101000011    0110011101000100    0110011101000101    0110011101000110    0110011101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26435 - 26439

  --0110011101001000    0110011101001001    0110011101001010    0110011101001011    0110011101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26440 - 26444

  --0110011101001101    0110011101001110    0110011101001111    0110011101010000    0110011101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26445 - 26449

  --0110011101010010    0110011101010011    0110011101010100    0110011101010101    0110011101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26450 - 26454

  --0110011101010111    0110011101011000    0110011101011001    0110011101011010    0110011101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26455 - 26459

  --0110011101011100    0110011101011101    0110011101011110    0110011101011111    0110011101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26460 - 26464

  --0110011101100001    0110011101100010    0110011101100011    0110011101100100    0110011101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26465 - 26469

  --0110011101100110    0110011101100111    0110011101101000    0110011101101001    0110011101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26470 - 26474

  --0110011101101011    0110011101101100    0110011101101101    0110011101101110    0110011101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26475 - 26479

  --0110011101110000    0110011101110001    0110011101110010    0110011101110011    0110011101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26480 - 26484

  --0110011101110101    0110011101110110    0110011101110111    0110011101111000    0110011101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26485 - 26489

  --0110011101111010    0110011101111011    0110011101111100    0110011101111101    0110011101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26490 - 26494

  --0110011101111111    0110011110000000    0110011110000001    0110011110000010    0110011110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26495 - 26499

  --0110011110000100    0110011110000101    0110011110000110    0110011110000111    0110011110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26500 - 26504

  --0110011110001001    0110011110001010    0110011110001011    0110011110001100    0110011110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26505 - 26509

  --0110011110001110    0110011110001111    0110011110010000    0110011110010001    0110011110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26510 - 26514

  --0110011110010011    0110011110010100    0110011110010101    0110011110010110    0110011110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26515 - 26519

  --0110011110011000    0110011110011001    0110011110011010    0110011110011011    0110011110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26520 - 26524

  --0110011110011101    0110011110011110    0110011110011111    0110011110100000    0110011110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26525 - 26529

  --0110011110100010    0110011110100011    0110011110100100    0110011110100101    0110011110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26530 - 26534

  --0110011110100111    0110011110101000    0110011110101001    0110011110101010    0110011110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26535 - 26539

  --0110011110101100    0110011110101101    0110011110101110    0110011110101111    0110011110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26540 - 26544

  --0110011110110001    0110011110110010    0110011110110011    0110011110110100    0110011110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26545 - 26549

  --0110011110110110    0110011110110111    0110011110111000    0110011110111001    0110011110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26550 - 26554

  --0110011110111011    0110011110111100    0110011110111101    0110011110111110    0110011110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26555 - 26559

  --0110011111000000    0110011111000001    0110011111000010    0110011111000011    0110011111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26560 - 26564

  --0110011111000101    0110011111000110    0110011111000111    0110011111001000    0110011111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26565 - 26569

  --0110011111001010    0110011111001011    0110011111001100    0110011111001101    0110011111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26570 - 26574

  --0110011111001111    0110011111010000    0110011111010001    0110011111010010    0110011111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26575 - 26579

  --0110011111010100    0110011111010101    0110011111010110    0110011111010111    0110011111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26580 - 26584

  --0110011111011001    0110011111011010    0110011111011011    0110011111011100    0110011111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26585 - 26589

  --0110011111011110    0110011111011111    0110011111100000    0110011111100001    0110011111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26590 - 26594

  --0110011111100011    0110011111100100    0110011111100101    0110011111100110    0110011111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26595 - 26599

  --0110011111101000    0110011111101001    0110011111101010    0110011111101011    0110011111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26600 - 26604

  --0110011111101101    0110011111101110    0110011111101111    0110011111110000    0110011111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26605 - 26609

  --0110011111110010    0110011111110011    0110011111110100    0110011111110101    0110011111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26610 - 26614

  --0110011111110111    0110011111111000    0110011111111001    0110011111111010    0110011111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26615 - 26619

  --0110011111111100    0110011111111101    0110011111111110    0110011111111111    0110100000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26620 - 26624

  --0110100000000001    0110100000000010    0110100000000011    0110100000000100    0110100000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26625 - 26629

  --0110100000000110    0110100000000111    0110100000001000    0110100000001001    0110100000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26630 - 26634

  --0110100000001011    0110100000001100    0110100000001101    0110100000001110    0110100000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26635 - 26639

  --0110100000010000    0110100000010001    0110100000010010    0110100000010011    0110100000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26640 - 26644

  --0110100000010101    0110100000010110    0110100000010111    0110100000011000    0110100000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26645 - 26649

  --0110100000011010    0110100000011011    0110100000011100    0110100000011101    0110100000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26650 - 26654

  --0110100000011111    0110100000100000    0110100000100001    0110100000100010    0110100000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26655 - 26659

  --0110100000100100    0110100000100101    0110100000100110    0110100000100111    0110100000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26660 - 26664

  --0110100000101001    0110100000101010    0110100000101011    0110100000101100    0110100000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26665 - 26669

  --0110100000101110    0110100000101111    0110100000110000    0110100000110001    0110100000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26670 - 26674

  --0110100000110011    0110100000110100    0110100000110101    0110100000110110    0110100000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26675 - 26679

  --0110100000111000    0110100000111001    0110100000111010    0110100000111011    0110100000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26680 - 26684

  --0110100000111101    0110100000111110    0110100000111111    0110100001000000    0110100001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26685 - 26689

  --0110100001000010    0110100001000011    0110100001000100    0110100001000101    0110100001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26690 - 26694

  --0110100001000111    0110100001001000    0110100001001001    0110100001001010    0110100001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26695 - 26699

  --0110100001001100    0110100001001101    0110100001001110    0110100001001111    0110100001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26700 - 26704

  --0110100001010001    0110100001010010    0110100001010011    0110100001010100    0110100001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26705 - 26709

  --0110100001010110    0110100001010111    0110100001011000    0110100001011001    0110100001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26710 - 26714

  --0110100001011011    0110100001011100    0110100001011101    0110100001011110    0110100001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26715 - 26719

  --0110100001100000    0110100001100001    0110100001100010    0110100001100011    0110100001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26720 - 26724

  --0110100001100101    0110100001100110    0110100001100111    0110100001101000    0110100001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26725 - 26729

  --0110100001101010    0110100001101011    0110100001101100    0110100001101101    0110100001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26730 - 26734

  --0110100001101111    0110100001110000    0110100001110001    0110100001110010    0110100001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26735 - 26739

  --0110100001110100    0110100001110101    0110100001110110    0110100001110111    0110100001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26740 - 26744

  --0110100001111001    0110100001111010    0110100001111011    0110100001111100    0110100001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26745 - 26749

  --0110100001111110    0110100001111111    0110100010000000    0110100010000001    0110100010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26750 - 26754

  --0110100010000011    0110100010000100    0110100010000101    0110100010000110    0110100010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26755 - 26759

  --0110100010001000    0110100010001001    0110100010001010    0110100010001011    0110100010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26760 - 26764

  --0110100010001101    0110100010001110    0110100010001111    0110100010010000    0110100010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26765 - 26769

  --0110100010010010    0110100010010011    0110100010010100    0110100010010101    0110100010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26770 - 26774

  --0110100010010111    0110100010011000    0110100010011001    0110100010011010    0110100010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26775 - 26779

  --0110100010011100    0110100010011101    0110100010011110    0110100010011111    0110100010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26780 - 26784

  --0110100010100001    0110100010100010    0110100010100011    0110100010100100    0110100010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26785 - 26789

  --0110100010100110    0110100010100111    0110100010101000    0110100010101001    0110100010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26790 - 26794

  --0110100010101011    0110100010101100    0110100010101101    0110100010101110    0110100010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26795 - 26799

  --0110100010110000    0110100010110001    0110100010110010    0110100010110011    0110100010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26800 - 26804

  --0110100010110101    0110100010110110    0110100010110111    0110100010111000    0110100010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26805 - 26809

  --0110100010111010    0110100010111011    0110100010111100    0110100010111101    0110100010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26810 - 26814

  --0110100010111111    0110100011000000    0110100011000001    0110100011000010    0110100011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26815 - 26819

  --0110100011000100    0110100011000101    0110100011000110    0110100011000111    0110100011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26820 - 26824

  --0110100011001001    0110100011001010    0110100011001011    0110100011001100    0110100011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26825 - 26829

  --0110100011001110    0110100011001111    0110100011010000    0110100011010001    0110100011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26830 - 26834

  --0110100011010011    0110100011010100    0110100011010101    0110100011010110    0110100011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26835 - 26839

  --0110100011011000    0110100011011001    0110100011011010    0110100011011011    0110100011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26840 - 26844

  --0110100011011101    0110100011011110    0110100011011111    0110100011100000    0110100011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26845 - 26849

  --0110100011100010    0110100011100011    0110100011100100    0110100011100101    0110100011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26850 - 26854

  --0110100011100111    0110100011101000    0110100011101001    0110100011101010    0110100011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26855 - 26859

  --0110100011101100    0110100011101101    0110100011101110    0110100011101111    0110100011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26860 - 26864

  --0110100011110001    0110100011110010    0110100011110011    0110100011110100    0110100011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26865 - 26869

  --0110100011110110    0110100011110111    0110100011111000    0110100011111001    0110100011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26870 - 26874

  --0110100011111011    0110100011111100    0110100011111101    0110100011111110    0110100011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26875 - 26879

  --0110100100000000    0110100100000001    0110100100000010    0110100100000011    0110100100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26880 - 26884

  --0110100100000101    0110100100000110    0110100100000111    0110100100001000    0110100100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26885 - 26889

  --0110100100001010    0110100100001011    0110100100001100    0110100100001101    0110100100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26890 - 26894

  --0110100100001111    0110100100010000    0110100100010001    0110100100010010    0110100100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26895 - 26899

  --0110100100010100    0110100100010101    0110100100010110    0110100100010111    0110100100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26900 - 26904

  --0110100100011001    0110100100011010    0110100100011011    0110100100011100    0110100100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26905 - 26909

  --0110100100011110    0110100100011111    0110100100100000    0110100100100001    0110100100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26910 - 26914

  --0110100100100011    0110100100100100    0110100100100101    0110100100100110    0110100100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26915 - 26919

  --0110100100101000    0110100100101001    0110100100101010    0110100100101011    0110100100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26920 - 26924

  --0110100100101101    0110100100101110    0110100100101111    0110100100110000    0110100100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26925 - 26929

  --0110100100110010    0110100100110011    0110100100110100    0110100100110101    0110100100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26930 - 26934

  --0110100100110111    0110100100111000    0110100100111001    0110100100111010    0110100100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26935 - 26939

  --0110100100111100    0110100100111101    0110100100111110    0110100100111111    0110100101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26940 - 26944

  --0110100101000001    0110100101000010    0110100101000011    0110100101000100    0110100101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26945 - 26949

  --0110100101000110    0110100101000111    0110100101001000    0110100101001001    0110100101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26950 - 26954

  --0110100101001011    0110100101001100    0110100101001101    0110100101001110    0110100101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26955 - 26959

  --0110100101010000    0110100101010001    0110100101010010    0110100101010011    0110100101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26960 - 26964

  --0110100101010101    0110100101010110    0110100101010111    0110100101011000    0110100101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26965 - 26969

  --0110100101011010    0110100101011011    0110100101011100    0110100101011101    0110100101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26970 - 26974

  --0110100101011111    0110100101100000    0110100101100001    0110100101100010    0110100101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26975 - 26979

  --0110100101100100    0110100101100101    0110100101100110    0110100101100111    0110100101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26980 - 26984

  --0110100101101001    0110100101101010    0110100101101011    0110100101101100    0110100101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26985 - 26989

  --0110100101101110    0110100101101111    0110100101110000    0110100101110001    0110100101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26990 - 26994

  --0110100101110011    0110100101110100    0110100101110101    0110100101110110    0110100101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 26995 - 26999

  --0110100101111000    0110100101111001    0110100101111010    0110100101111011    0110100101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27000 - 27004

  --0110100101111101    0110100101111110    0110100101111111    0110100110000000    0110100110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27005 - 27009

  --0110100110000010    0110100110000011    0110100110000100    0110100110000101    0110100110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27010 - 27014

  --0110100110000111    0110100110001000    0110100110001001    0110100110001010    0110100110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27015 - 27019

  --0110100110001100    0110100110001101    0110100110001110    0110100110001111    0110100110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27020 - 27024

  --0110100110010001    0110100110010010    0110100110010011    0110100110010100    0110100110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27025 - 27029

  --0110100110010110    0110100110010111    0110100110011000    0110100110011001    0110100110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27030 - 27034

  --0110100110011011    0110100110011100    0110100110011101    0110100110011110    0110100110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27035 - 27039

  --0110100110100000    0110100110100001    0110100110100010    0110100110100011    0110100110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27040 - 27044

  --0110100110100101    0110100110100110    0110100110100111    0110100110101000    0110100110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27045 - 27049

  --0110100110101010    0110100110101011    0110100110101100    0110100110101101    0110100110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27050 - 27054

  --0110100110101111    0110100110110000    0110100110110001    0110100110110010    0110100110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27055 - 27059

  --0110100110110100    0110100110110101    0110100110110110    0110100110110111    0110100110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27060 - 27064

  --0110100110111001    0110100110111010    0110100110111011    0110100110111100    0110100110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27065 - 27069

  --0110100110111110    0110100110111111    0110100111000000    0110100111000001    0110100111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27070 - 27074

  --0110100111000011    0110100111000100    0110100111000101    0110100111000110    0110100111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27075 - 27079

  --0110100111001000    0110100111001001    0110100111001010    0110100111001011    0110100111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27080 - 27084

  --0110100111001101    0110100111001110    0110100111001111    0110100111010000    0110100111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27085 - 27089

  --0110100111010010    0110100111010011    0110100111010100    0110100111010101    0110100111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27090 - 27094

  --0110100111010111    0110100111011000    0110100111011001    0110100111011010    0110100111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27095 - 27099

  --0110100111011100    0110100111011101    0110100111011110    0110100111011111    0110100111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27100 - 27104

  --0110100111100001    0110100111100010    0110100111100011    0110100111100100    0110100111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27105 - 27109

  --0110100111100110    0110100111100111    0110100111101000    0110100111101001    0110100111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27110 - 27114

  --0110100111101011    0110100111101100    0110100111101101    0110100111101110    0110100111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27115 - 27119

  --0110100111110000    0110100111110001    0110100111110010    0110100111110011    0110100111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27120 - 27124

  --0110100111110101    0110100111110110    0110100111110111    0110100111111000    0110100111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27125 - 27129

  --0110100111111010    0110100111111011    0110100111111100    0110100111111101    0110100111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27130 - 27134

  --0110100111111111    0110101000000000    0110101000000001    0110101000000010    0110101000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27135 - 27139

  --0110101000000100    0110101000000101    0110101000000110    0110101000000111    0110101000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27140 - 27144

  --0110101000001001    0110101000001010    0110101000001011    0110101000001100    0110101000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27145 - 27149

  --0110101000001110    0110101000001111    0110101000010000    0110101000010001    0110101000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27150 - 27154

  --0110101000010011    0110101000010100    0110101000010101    0110101000010110    0110101000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27155 - 27159

  --0110101000011000    0110101000011001    0110101000011010    0110101000011011    0110101000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27160 - 27164

  --0110101000011101    0110101000011110    0110101000011111    0110101000100000    0110101000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27165 - 27169

  --0110101000100010    0110101000100011    0110101000100100    0110101000100101    0110101000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27170 - 27174

  --0110101000100111    0110101000101000    0110101000101001    0110101000101010    0110101000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27175 - 27179

  --0110101000101100    0110101000101101    0110101000101110    0110101000101111    0110101000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27180 - 27184

  --0110101000110001    0110101000110010    0110101000110011    0110101000110100    0110101000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27185 - 27189

  --0110101000110110    0110101000110111    0110101000111000    0110101000111001    0110101000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27190 - 27194

  --0110101000111011    0110101000111100    0110101000111101    0110101000111110    0110101000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27195 - 27199

  --0110101001000000    0110101001000001    0110101001000010    0110101001000011    0110101001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27200 - 27204

  --0110101001000101    0110101001000110    0110101001000111    0110101001001000    0110101001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27205 - 27209

  --0110101001001010    0110101001001011    0110101001001100    0110101001001101    0110101001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27210 - 27214

  --0110101001001111    0110101001010000    0110101001010001    0110101001010010    0110101001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27215 - 27219

  --0110101001010100    0110101001010101    0110101001010110    0110101001010111    0110101001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27220 - 27224

  --0110101001011001    0110101001011010    0110101001011011    0110101001011100    0110101001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27225 - 27229

  --0110101001011110    0110101001011111    0110101001100000    0110101001100001    0110101001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27230 - 27234

  --0110101001100011    0110101001100100    0110101001100101    0110101001100110    0110101001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27235 - 27239

  --0110101001101000    0110101001101001    0110101001101010    0110101001101011    0110101001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27240 - 27244

  --0110101001101101    0110101001101110    0110101001101111    0110101001110000    0110101001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27245 - 27249

  --0110101001110010    0110101001110011    0110101001110100    0110101001110101    0110101001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27250 - 27254

  --0110101001110111    0110101001111000    0110101001111001    0110101001111010    0110101001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27255 - 27259

  --0110101001111100    0110101001111101    0110101001111110    0110101001111111    0110101010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27260 - 27264

  --0110101010000001    0110101010000010    0110101010000011    0110101010000100    0110101010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27265 - 27269

  --0110101010000110    0110101010000111    0110101010001000    0110101010001001    0110101010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27270 - 27274

  --0110101010001011    0110101010001100    0110101010001101    0110101010001110    0110101010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27275 - 27279

  --0110101010010000    0110101010010001    0110101010010010    0110101010010011    0110101010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27280 - 27284

  --0110101010010101    0110101010010110    0110101010010111    0110101010011000    0110101010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27285 - 27289

  --0110101010011010    0110101010011011    0110101010011100    0110101010011101    0110101010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27290 - 27294

  --0110101010011111    0110101010100000    0110101010100001    0110101010100010    0110101010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27295 - 27299

  --0110101010100100    0110101010100101    0110101010100110    0110101010100111    0110101010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27300 - 27304

  --0110101010101001    0110101010101010    0110101010101011    0110101010101100    0110101010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27305 - 27309

  --0110101010101110    0110101010101111    0110101010110000    0110101010110001    0110101010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27310 - 27314

  --0110101010110011    0110101010110100    0110101010110101    0110101010110110    0110101010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27315 - 27319

  --0110101010111000    0110101010111001    0110101010111010    0110101010111011    0110101010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27320 - 27324

  --0110101010111101    0110101010111110    0110101010111111    0110101011000000    0110101011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27325 - 27329

  --0110101011000010    0110101011000011    0110101011000100    0110101011000101    0110101011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27330 - 27334

  --0110101011000111    0110101011001000    0110101011001001    0110101011001010    0110101011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27335 - 27339

  --0110101011001100    0110101011001101    0110101011001110    0110101011001111    0110101011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27340 - 27344

  --0110101011010001    0110101011010010    0110101011010011    0110101011010100    0110101011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27345 - 27349

  --0110101011010110    0110101011010111    0110101011011000    0110101011011001    0110101011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27350 - 27354

  --0110101011011011    0110101011011100    0110101011011101    0110101011011110    0110101011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27355 - 27359

  --0110101011100000    0110101011100001    0110101011100010    0110101011100011    0110101011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27360 - 27364

  --0110101011100101    0110101011100110    0110101011100111    0110101011101000    0110101011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27365 - 27369

  --0110101011101010    0110101011101011    0110101011101100    0110101011101101    0110101011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27370 - 27374

  --0110101011101111    0110101011110000    0110101011110001    0110101011110010    0110101011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27375 - 27379

  --0110101011110100    0110101011110101    0110101011110110    0110101011110111    0110101011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27380 - 27384

  --0110101011111001    0110101011111010    0110101011111011    0110101011111100    0110101011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27385 - 27389

  --0110101011111110    0110101011111111    0110101100000000    0110101100000001    0110101100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27390 - 27394

  --0110101100000011    0110101100000100    0110101100000101    0110101100000110    0110101100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27395 - 27399

  --0110101100001000    0110101100001001    0110101100001010    0110101100001011    0110101100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27400 - 27404

  --0110101100001101    0110101100001110    0110101100001111    0110101100010000    0110101100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27405 - 27409

  --0110101100010010    0110101100010011    0110101100010100    0110101100010101    0110101100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27410 - 27414

  --0110101100010111    0110101100011000    0110101100011001    0110101100011010    0110101100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27415 - 27419

  --0110101100011100    0110101100011101    0110101100011110    0110101100011111    0110101100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27420 - 27424

  --0110101100100001    0110101100100010    0110101100100011    0110101100100100    0110101100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27425 - 27429

  --0110101100100110    0110101100100111    0110101100101000    0110101100101001    0110101100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27430 - 27434

  --0110101100101011    0110101100101100    0110101100101101    0110101100101110    0110101100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27435 - 27439

  --0110101100110000    0110101100110001    0110101100110010    0110101100110011    0110101100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27440 - 27444

  --0110101100110101    0110101100110110    0110101100110111    0110101100111000    0110101100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27445 - 27449

  --0110101100111010    0110101100111011    0110101100111100    0110101100111101    0110101100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27450 - 27454

  --0110101100111111    0110101101000000    0110101101000001    0110101101000010    0110101101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27455 - 27459

  --0110101101000100    0110101101000101    0110101101000110    0110101101000111    0110101101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27460 - 27464

  --0110101101001001    0110101101001010    0110101101001011    0110101101001100    0110101101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27465 - 27469

  --0110101101001110    0110101101001111    0110101101010000    0110101101010001    0110101101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27470 - 27474

  --0110101101010011    0110101101010100    0110101101010101    0110101101010110    0110101101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27475 - 27479

  --0110101101011000    0110101101011001    0110101101011010    0110101101011011    0110101101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27480 - 27484

  --0110101101011101    0110101101011110    0110101101011111    0110101101100000    0110101101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27485 - 27489

  --0110101101100010    0110101101100011    0110101101100100    0110101101100101    0110101101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27490 - 27494

  --0110101101100111    0110101101101000    0110101101101001    0110101101101010    0110101101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27495 - 27499

  --0110101101101100    0110101101101101    0110101101101110    0110101101101111    0110101101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27500 - 27504

  --0110101101110001    0110101101110010    0110101101110011    0110101101110100    0110101101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27505 - 27509

  --0110101101110110    0110101101110111    0110101101111000    0110101101111001    0110101101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27510 - 27514

  --0110101101111011    0110101101111100    0110101101111101    0110101101111110    0110101101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27515 - 27519

  --0110101110000000    0110101110000001    0110101110000010    0110101110000011    0110101110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27520 - 27524

  --0110101110000101    0110101110000110    0110101110000111    0110101110001000    0110101110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27525 - 27529

  --0110101110001010    0110101110001011    0110101110001100    0110101110001101    0110101110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27530 - 27534

  --0110101110001111    0110101110010000    0110101110010001    0110101110010010    0110101110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27535 - 27539

  --0110101110010100    0110101110010101    0110101110010110    0110101110010111    0110101110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27540 - 27544

  --0110101110011001    0110101110011010    0110101110011011    0110101110011100    0110101110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27545 - 27549

  --0110101110011110    0110101110011111    0110101110100000    0110101110100001    0110101110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27550 - 27554

  --0110101110100011    0110101110100100    0110101110100101    0110101110100110    0110101110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27555 - 27559

  --0110101110101000    0110101110101001    0110101110101010    0110101110101011    0110101110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27560 - 27564

  --0110101110101101    0110101110101110    0110101110101111    0110101110110000    0110101110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27565 - 27569

  --0110101110110010    0110101110110011    0110101110110100    0110101110110101    0110101110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27570 - 27574

  --0110101110110111    0110101110111000    0110101110111001    0110101110111010    0110101110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27575 - 27579

  --0110101110111100    0110101110111101    0110101110111110    0110101110111111    0110101111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27580 - 27584

  --0110101111000001    0110101111000010    0110101111000011    0110101111000100    0110101111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27585 - 27589

  --0110101111000110    0110101111000111    0110101111001000    0110101111001001    0110101111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27590 - 27594

  --0110101111001011    0110101111001100    0110101111001101    0110101111001110    0110101111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27595 - 27599

  --0110101111010000    0110101111010001    0110101111010010    0110101111010011    0110101111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27600 - 27604

  --0110101111010101    0110101111010110    0110101111010111    0110101111011000    0110101111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27605 - 27609

  --0110101111011010    0110101111011011    0110101111011100    0110101111011101    0110101111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27610 - 27614

  --0110101111011111    0110101111100000    0110101111100001    0110101111100010    0110101111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27615 - 27619

  --0110101111100100    0110101111100101    0110101111100110    0110101111100111    0110101111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27620 - 27624

  --0110101111101001    0110101111101010    0110101111101011    0110101111101100    0110101111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27625 - 27629

  --0110101111101110    0110101111101111    0110101111110000    0110101111110001    0110101111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27630 - 27634

  --0110101111110011    0110101111110100    0110101111110101    0110101111110110    0110101111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27635 - 27639

  --0110101111111000    0110101111111001    0110101111111010    0110101111111011    0110101111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27640 - 27644

  --0110101111111101    0110101111111110    0110101111111111    0110110000000000    0110110000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27645 - 27649

  --0110110000000010    0110110000000011    0110110000000100    0110110000000101    0110110000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27650 - 27654

  --0110110000000111    0110110000001000    0110110000001001    0110110000001010    0110110000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27655 - 27659

  --0110110000001100    0110110000001101    0110110000001110    0110110000001111    0110110000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27660 - 27664

  --0110110000010001    0110110000010010    0110110000010011    0110110000010100    0110110000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27665 - 27669

  --0110110000010110    0110110000010111    0110110000011000    0110110000011001    0110110000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27670 - 27674

  --0110110000011011    0110110000011100    0110110000011101    0110110000011110    0110110000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27675 - 27679

  --0110110000100000    0110110000100001    0110110000100010    0110110000100011    0110110000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27680 - 27684

  --0110110000100101    0110110000100110    0110110000100111    0110110000101000    0110110000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27685 - 27689

  --0110110000101010    0110110000101011    0110110000101100    0110110000101101    0110110000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27690 - 27694

  --0110110000101111    0110110000110000    0110110000110001    0110110000110010    0110110000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27695 - 27699

  --0110110000110100    0110110000110101    0110110000110110    0110110000110111    0110110000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27700 - 27704

  --0110110000111001    0110110000111010    0110110000111011    0110110000111100    0110110000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27705 - 27709

  --0110110000111110    0110110000111111    0110110001000000    0110110001000001    0110110001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27710 - 27714

  --0110110001000011    0110110001000100    0110110001000101    0110110001000110    0110110001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27715 - 27719

  --0110110001001000    0110110001001001    0110110001001010    0110110001001011    0110110001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27720 - 27724

  --0110110001001101    0110110001001110    0110110001001111    0110110001010000    0110110001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27725 - 27729

  --0110110001010010    0110110001010011    0110110001010100    0110110001010101    0110110001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27730 - 27734

  --0110110001010111    0110110001011000    0110110001011001    0110110001011010    0110110001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27735 - 27739

  --0110110001011100    0110110001011101    0110110001011110    0110110001011111    0110110001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27740 - 27744

  --0110110001100001    0110110001100010    0110110001100011    0110110001100100    0110110001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27745 - 27749

  --0110110001100110    0110110001100111    0110110001101000    0110110001101001    0110110001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27750 - 27754

  --0110110001101011    0110110001101100    0110110001101101    0110110001101110    0110110001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27755 - 27759

  --0110110001110000    0110110001110001    0110110001110010    0110110001110011    0110110001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27760 - 27764

  --0110110001110101    0110110001110110    0110110001110111    0110110001111000    0110110001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27765 - 27769

  --0110110001111010    0110110001111011    0110110001111100    0110110001111101    0110110001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27770 - 27774

  --0110110001111111    0110110010000000    0110110010000001    0110110010000010    0110110010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27775 - 27779

  --0110110010000100    0110110010000101    0110110010000110    0110110010000111    0110110010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27780 - 27784

  --0110110010001001    0110110010001010    0110110010001011    0110110010001100    0110110010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27785 - 27789

  --0110110010001110    0110110010001111    0110110010010000    0110110010010001    0110110010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27790 - 27794

  --0110110010010011    0110110010010100    0110110010010101    0110110010010110    0110110010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27795 - 27799

  --0110110010011000    0110110010011001    0110110010011010    0110110010011011    0110110010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27800 - 27804

  --0110110010011101    0110110010011110    0110110010011111    0110110010100000    0110110010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27805 - 27809

  --0110110010100010    0110110010100011    0110110010100100    0110110010100101    0110110010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27810 - 27814

  --0110110010100111    0110110010101000    0110110010101001    0110110010101010    0110110010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27815 - 27819

  --0110110010101100    0110110010101101    0110110010101110    0110110010101111    0110110010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27820 - 27824

  --0110110010110001    0110110010110010    0110110010110011    0110110010110100    0110110010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27825 - 27829

  --0110110010110110    0110110010110111    0110110010111000    0110110010111001    0110110010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27830 - 27834

  --0110110010111011    0110110010111100    0110110010111101    0110110010111110    0110110010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27835 - 27839

  --0110110011000000    0110110011000001    0110110011000010    0110110011000011    0110110011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27840 - 27844

  --0110110011000101    0110110011000110    0110110011000111    0110110011001000    0110110011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27845 - 27849

  --0110110011001010    0110110011001011    0110110011001100    0110110011001101    0110110011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27850 - 27854

  --0110110011001111    0110110011010000    0110110011010001    0110110011010010    0110110011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27855 - 27859

  --0110110011010100    0110110011010101    0110110011010110    0110110011010111    0110110011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27860 - 27864

  --0110110011011001    0110110011011010    0110110011011011    0110110011011100    0110110011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27865 - 27869

  --0110110011011110    0110110011011111    0110110011100000    0110110011100001    0110110011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27870 - 27874

  --0110110011100011    0110110011100100    0110110011100101    0110110011100110    0110110011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27875 - 27879

  --0110110011101000    0110110011101001    0110110011101010    0110110011101011    0110110011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27880 - 27884

  --0110110011101101    0110110011101110    0110110011101111    0110110011110000    0110110011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27885 - 27889

  --0110110011110010    0110110011110011    0110110011110100    0110110011110101    0110110011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27890 - 27894

  --0110110011110111    0110110011111000    0110110011111001    0110110011111010    0110110011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27895 - 27899

  --0110110011111100    0110110011111101    0110110011111110    0110110011111111    0110110100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27900 - 27904

  --0110110100000001    0110110100000010    0110110100000011    0110110100000100    0110110100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27905 - 27909

  --0110110100000110    0110110100000111    0110110100001000    0110110100001001    0110110100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27910 - 27914

  --0110110100001011    0110110100001100    0110110100001101    0110110100001110    0110110100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27915 - 27919

  --0110110100010000    0110110100010001    0110110100010010    0110110100010011    0110110100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27920 - 27924

  --0110110100010101    0110110100010110    0110110100010111    0110110100011000    0110110100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27925 - 27929

  --0110110100011010    0110110100011011    0110110100011100    0110110100011101    0110110100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27930 - 27934

  --0110110100011111    0110110100100000    0110110100100001    0110110100100010    0110110100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27935 - 27939

  --0110110100100100    0110110100100101    0110110100100110    0110110100100111    0110110100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27940 - 27944

  --0110110100101001    0110110100101010    0110110100101011    0110110100101100    0110110100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27945 - 27949

  --0110110100101110    0110110100101111    0110110100110000    0110110100110001    0110110100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27950 - 27954

  --0110110100110011    0110110100110100    0110110100110101    0110110100110110    0110110100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27955 - 27959

  --0110110100111000    0110110100111001    0110110100111010    0110110100111011    0110110100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27960 - 27964

  --0110110100111101    0110110100111110    0110110100111111    0110110101000000    0110110101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27965 - 27969

  --0110110101000010    0110110101000011    0110110101000100    0110110101000101    0110110101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27970 - 27974

  --0110110101000111    0110110101001000    0110110101001001    0110110101001010    0110110101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27975 - 27979

  --0110110101001100    0110110101001101    0110110101001110    0110110101001111    0110110101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27980 - 27984

  --0110110101010001    0110110101010010    0110110101010011    0110110101010100    0110110101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27985 - 27989

  --0110110101010110    0110110101010111    0110110101011000    0110110101011001    0110110101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27990 - 27994

  --0110110101011011    0110110101011100    0110110101011101    0110110101011110    0110110101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 27995 - 27999

  --0110110101100000    0110110101100001    0110110101100010    0110110101100011    0110110101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28000 - 28004

  --0110110101100101    0110110101100110    0110110101100111    0110110101101000    0110110101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28005 - 28009

  --0110110101101010    0110110101101011    0110110101101100    0110110101101101    0110110101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28010 - 28014

  --0110110101101111    0110110101110000    0110110101110001    0110110101110010    0110110101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28015 - 28019

  --0110110101110100    0110110101110101    0110110101110110    0110110101110111    0110110101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28020 - 28024

  --0110110101111001    0110110101111010    0110110101111011    0110110101111100    0110110101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28025 - 28029

  --0110110101111110    0110110101111111    0110110110000000    0110110110000001    0110110110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28030 - 28034

  --0110110110000011    0110110110000100    0110110110000101    0110110110000110    0110110110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28035 - 28039

  --0110110110001000    0110110110001001    0110110110001010    0110110110001011    0110110110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28040 - 28044

  --0110110110001101    0110110110001110    0110110110001111    0110110110010000    0110110110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28045 - 28049

  --0110110110010010    0110110110010011    0110110110010100    0110110110010101    0110110110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28050 - 28054

  --0110110110010111    0110110110011000    0110110110011001    0110110110011010    0110110110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28055 - 28059

  --0110110110011100    0110110110011101    0110110110011110    0110110110011111    0110110110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28060 - 28064

  --0110110110100001    0110110110100010    0110110110100011    0110110110100100    0110110110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28065 - 28069

  --0110110110100110    0110110110100111    0110110110101000    0110110110101001    0110110110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28070 - 28074

  --0110110110101011    0110110110101100    0110110110101101    0110110110101110    0110110110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28075 - 28079

  --0110110110110000    0110110110110001    0110110110110010    0110110110110011    0110110110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28080 - 28084

  --0110110110110101    0110110110110110    0110110110110111    0110110110111000    0110110110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28085 - 28089

  --0110110110111010    0110110110111011    0110110110111100    0110110110111101    0110110110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28090 - 28094

  --0110110110111111    0110110111000000    0110110111000001    0110110111000010    0110110111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28095 - 28099

  --0110110111000100    0110110111000101    0110110111000110    0110110111000111    0110110111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28100 - 28104

  --0110110111001001    0110110111001010    0110110111001011    0110110111001100    0110110111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28105 - 28109

  --0110110111001110    0110110111001111    0110110111010000    0110110111010001    0110110111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28110 - 28114

  --0110110111010011    0110110111010100    0110110111010101    0110110111010110    0110110111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28115 - 28119

  --0110110111011000    0110110111011001    0110110111011010    0110110111011011    0110110111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28120 - 28124

  --0110110111011101    0110110111011110    0110110111011111    0110110111100000    0110110111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28125 - 28129

  --0110110111100010    0110110111100011    0110110111100100    0110110111100101    0110110111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28130 - 28134

  --0110110111100111    0110110111101000    0110110111101001    0110110111101010    0110110111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28135 - 28139

  --0110110111101100    0110110111101101    0110110111101110    0110110111101111    0110110111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28140 - 28144

  --0110110111110001    0110110111110010    0110110111110011    0110110111110100    0110110111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28145 - 28149

  --0110110111110110    0110110111110111    0110110111111000    0110110111111001    0110110111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28150 - 28154

  --0110110111111011    0110110111111100    0110110111111101    0110110111111110    0110110111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28155 - 28159

  --0110111000000000    0110111000000001    0110111000000010    0110111000000011    0110111000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28160 - 28164

  --0110111000000101    0110111000000110    0110111000000111    0110111000001000    0110111000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28165 - 28169

  --0110111000001010    0110111000001011    0110111000001100    0110111000001101    0110111000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28170 - 28174

  --0110111000001111    0110111000010000    0110111000010001    0110111000010010    0110111000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28175 - 28179

  --0110111000010100    0110111000010101    0110111000010110    0110111000010111    0110111000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28180 - 28184

  --0110111000011001    0110111000011010    0110111000011011    0110111000011100    0110111000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28185 - 28189

  --0110111000011110    0110111000011111    0110111000100000    0110111000100001    0110111000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28190 - 28194

  --0110111000100011    0110111000100100    0110111000100101    0110111000100110    0110111000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28195 - 28199

  --0110111000101000    0110111000101001    0110111000101010    0110111000101011    0110111000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28200 - 28204

  --0110111000101101    0110111000101110    0110111000101111    0110111000110000    0110111000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28205 - 28209

  --0110111000110010    0110111000110011    0110111000110100    0110111000110101    0110111000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28210 - 28214

  --0110111000110111    0110111000111000    0110111000111001    0110111000111010    0110111000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28215 - 28219

  --0110111000111100    0110111000111101    0110111000111110    0110111000111111    0110111001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28220 - 28224

  --0110111001000001    0110111001000010    0110111001000011    0110111001000100    0110111001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28225 - 28229

  --0110111001000110    0110111001000111    0110111001001000    0110111001001001    0110111001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28230 - 28234

  --0110111001001011    0110111001001100    0110111001001101    0110111001001110    0110111001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28235 - 28239

  --0110111001010000    0110111001010001    0110111001010010    0110111001010011    0110111001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28240 - 28244

  --0110111001010101    0110111001010110    0110111001010111    0110111001011000    0110111001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28245 - 28249

  --0110111001011010    0110111001011011    0110111001011100    0110111001011101    0110111001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28250 - 28254

  --0110111001011111    0110111001100000    0110111001100001    0110111001100010    0110111001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28255 - 28259

  --0110111001100100    0110111001100101    0110111001100110    0110111001100111    0110111001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28260 - 28264

  --0110111001101001    0110111001101010    0110111001101011    0110111001101100    0110111001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28265 - 28269

  --0110111001101110    0110111001101111    0110111001110000    0110111001110001    0110111001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28270 - 28274

  --0110111001110011    0110111001110100    0110111001110101    0110111001110110    0110111001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28275 - 28279

  --0110111001111000    0110111001111001    0110111001111010    0110111001111011    0110111001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28280 - 28284

  --0110111001111101    0110111001111110    0110111001111111    0110111010000000    0110111010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28285 - 28289

  --0110111010000010    0110111010000011    0110111010000100    0110111010000101    0110111010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28290 - 28294

  --0110111010000111    0110111010001000    0110111010001001    0110111010001010    0110111010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28295 - 28299

  --0110111010001100    0110111010001101    0110111010001110    0110111010001111    0110111010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28300 - 28304

  --0110111010010001    0110111010010010    0110111010010011    0110111010010100    0110111010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28305 - 28309

  --0110111010010110    0110111010010111    0110111010011000    0110111010011001    0110111010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28310 - 28314

  --0110111010011011    0110111010011100    0110111010011101    0110111010011110    0110111010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28315 - 28319

  --0110111010100000    0110111010100001    0110111010100010    0110111010100011    0110111010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28320 - 28324

  --0110111010100101    0110111010100110    0110111010100111    0110111010101000    0110111010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28325 - 28329

  --0110111010101010    0110111010101011    0110111010101100    0110111010101101    0110111010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28330 - 28334

  --0110111010101111    0110111010110000    0110111010110001    0110111010110010    0110111010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28335 - 28339

  --0110111010110100    0110111010110101    0110111010110110    0110111010110111    0110111010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28340 - 28344

  --0110111010111001    0110111010111010    0110111010111011    0110111010111100    0110111010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28345 - 28349

  --0110111010111110    0110111010111111    0110111011000000    0110111011000001    0110111011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28350 - 28354

  --0110111011000011    0110111011000100    0110111011000101    0110111011000110    0110111011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28355 - 28359

  --0110111011001000    0110111011001001    0110111011001010    0110111011001011    0110111011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28360 - 28364

  --0110111011001101    0110111011001110    0110111011001111    0110111011010000    0110111011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28365 - 28369

  --0110111011010010    0110111011010011    0110111011010100    0110111011010101    0110111011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28370 - 28374

  --0110111011010111    0110111011011000    0110111011011001    0110111011011010    0110111011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28375 - 28379

  --0110111011011100    0110111011011101    0110111011011110    0110111011011111    0110111011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28380 - 28384

  --0110111011100001    0110111011100010    0110111011100011    0110111011100100    0110111011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28385 - 28389

  --0110111011100110    0110111011100111    0110111011101000    0110111011101001    0110111011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28390 - 28394

  --0110111011101011    0110111011101100    0110111011101101    0110111011101110    0110111011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28395 - 28399

  --0110111011110000    0110111011110001    0110111011110010    0110111011110011    0110111011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28400 - 28404

  --0110111011110101    0110111011110110    0110111011110111    0110111011111000    0110111011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28405 - 28409

  --0110111011111010    0110111011111011    0110111011111100    0110111011111101    0110111011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28410 - 28414

  --0110111011111111    0110111100000000    0110111100000001    0110111100000010    0110111100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28415 - 28419

  --0110111100000100    0110111100000101    0110111100000110    0110111100000111    0110111100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28420 - 28424

  --0110111100001001    0110111100001010    0110111100001011    0110111100001100    0110111100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28425 - 28429

  --0110111100001110    0110111100001111    0110111100010000    0110111100010001    0110111100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28430 - 28434

  --0110111100010011    0110111100010100    0110111100010101    0110111100010110    0110111100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28435 - 28439

  --0110111100011000    0110111100011001    0110111100011010    0110111100011011    0110111100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28440 - 28444

  --0110111100011101    0110111100011110    0110111100011111    0110111100100000    0110111100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28445 - 28449

  --0110111100100010    0110111100100011    0110111100100100    0110111100100101    0110111100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28450 - 28454

  --0110111100100111    0110111100101000    0110111100101001    0110111100101010    0110111100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28455 - 28459

  --0110111100101100    0110111100101101    0110111100101110    0110111100101111    0110111100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28460 - 28464

  --0110111100110001    0110111100110010    0110111100110011    0110111100110100    0110111100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28465 - 28469

  --0110111100110110    0110111100110111    0110111100111000    0110111100111001    0110111100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28470 - 28474

  --0110111100111011    0110111100111100    0110111100111101    0110111100111110    0110111100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28475 - 28479

  --0110111101000000    0110111101000001    0110111101000010    0110111101000011    0110111101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28480 - 28484

  --0110111101000101    0110111101000110    0110111101000111    0110111101001000    0110111101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28485 - 28489

  --0110111101001010    0110111101001011    0110111101001100    0110111101001101    0110111101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28490 - 28494

  --0110111101001111    0110111101010000    0110111101010001    0110111101010010    0110111101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28495 - 28499

  --0110111101010100    0110111101010101    0110111101010110    0110111101010111    0110111101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28500 - 28504

  --0110111101011001    0110111101011010    0110111101011011    0110111101011100    0110111101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28505 - 28509

  --0110111101011110    0110111101011111    0110111101100000    0110111101100001    0110111101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28510 - 28514

  --0110111101100011    0110111101100100    0110111101100101    0110111101100110    0110111101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28515 - 28519

  --0110111101101000    0110111101101001    0110111101101010    0110111101101011    0110111101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28520 - 28524

  --0110111101101101    0110111101101110    0110111101101111    0110111101110000    0110111101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28525 - 28529

  --0110111101110010    0110111101110011    0110111101110100    0110111101110101    0110111101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28530 - 28534

  --0110111101110111    0110111101111000    0110111101111001    0110111101111010    0110111101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28535 - 28539

  --0110111101111100    0110111101111101    0110111101111110    0110111101111111    0110111110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28540 - 28544

  --0110111110000001    0110111110000010    0110111110000011    0110111110000100    0110111110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28545 - 28549

  --0110111110000110    0110111110000111    0110111110001000    0110111110001001    0110111110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28550 - 28554

  --0110111110001011    0110111110001100    0110111110001101    0110111110001110    0110111110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28555 - 28559

  --0110111110010000    0110111110010001    0110111110010010    0110111110010011    0110111110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28560 - 28564

  --0110111110010101    0110111110010110    0110111110010111    0110111110011000    0110111110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28565 - 28569

  --0110111110011010    0110111110011011    0110111110011100    0110111110011101    0110111110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28570 - 28574

  --0110111110011111    0110111110100000    0110111110100001    0110111110100010    0110111110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28575 - 28579

  --0110111110100100    0110111110100101    0110111110100110    0110111110100111    0110111110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28580 - 28584

  --0110111110101001    0110111110101010    0110111110101011    0110111110101100    0110111110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28585 - 28589

  --0110111110101110    0110111110101111    0110111110110000    0110111110110001    0110111110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28590 - 28594

  --0110111110110011    0110111110110100    0110111110110101    0110111110110110    0110111110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28595 - 28599

  --0110111110111000    0110111110111001    0110111110111010    0110111110111011    0110111110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28600 - 28604

  --0110111110111101    0110111110111110    0110111110111111    0110111111000000    0110111111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28605 - 28609

  --0110111111000010    0110111111000011    0110111111000100    0110111111000101    0110111111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28610 - 28614

  --0110111111000111    0110111111001000    0110111111001001    0110111111001010    0110111111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28615 - 28619

  --0110111111001100    0110111111001101    0110111111001110    0110111111001111    0110111111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28620 - 28624

  --0110111111010001    0110111111010010    0110111111010011    0110111111010100    0110111111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28625 - 28629

  --0110111111010110    0110111111010111    0110111111011000    0110111111011001    0110111111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28630 - 28634

  --0110111111011011    0110111111011100    0110111111011101    0110111111011110    0110111111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28635 - 28639

  --0110111111100000    0110111111100001    0110111111100010    0110111111100011    0110111111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28640 - 28644

  --0110111111100101    0110111111100110    0110111111100111    0110111111101000    0110111111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28645 - 28649

  --0110111111101010    0110111111101011    0110111111101100    0110111111101101    0110111111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28650 - 28654

  --0110111111101111    0110111111110000    0110111111110001    0110111111110010    0110111111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28655 - 28659

  --0110111111110100    0110111111110101    0110111111110110    0110111111110111    0110111111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28660 - 28664

  --0110111111111001    0110111111111010    0110111111111011    0110111111111100    0110111111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28665 - 28669

  --0110111111111110    0110111111111111    0111000000000000    0111000000000001    0111000000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28670 - 28674

  --0111000000000011    0111000000000100    0111000000000101    0111000000000110    0111000000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28675 - 28679

  --0111000000001000    0111000000001001    0111000000001010    0111000000001011    0111000000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28680 - 28684

  --0111000000001101    0111000000001110    0111000000001111    0111000000010000    0111000000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28685 - 28689

  --0111000000010010    0111000000010011    0111000000010100    0111000000010101    0111000000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28690 - 28694

  --0111000000010111    0111000000011000    0111000000011001    0111000000011010    0111000000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28695 - 28699

  --0111000000011100    0111000000011101    0111000000011110    0111000000011111    0111000000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28700 - 28704

  --0111000000100001    0111000000100010    0111000000100011    0111000000100100    0111000000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28705 - 28709

  --0111000000100110    0111000000100111    0111000000101000    0111000000101001    0111000000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28710 - 28714

  --0111000000101011    0111000000101100    0111000000101101    0111000000101110    0111000000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28715 - 28719

  --0111000000110000    0111000000110001    0111000000110010    0111000000110011    0111000000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28720 - 28724

  --0111000000110101    0111000000110110    0111000000110111    0111000000111000    0111000000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28725 - 28729

  --0111000000111010    0111000000111011    0111000000111100    0111000000111101    0111000000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28730 - 28734

  --0111000000111111    0111000001000000    0111000001000001    0111000001000010    0111000001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28735 - 28739

  --0111000001000100    0111000001000101    0111000001000110    0111000001000111    0111000001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28740 - 28744

  --0111000001001001    0111000001001010    0111000001001011    0111000001001100    0111000001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28745 - 28749

  --0111000001001110    0111000001001111    0111000001010000    0111000001010001    0111000001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28750 - 28754

  --0111000001010011    0111000001010100    0111000001010101    0111000001010110    0111000001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28755 - 28759

  --0111000001011000    0111000001011001    0111000001011010    0111000001011011    0111000001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28760 - 28764

  --0111000001011101    0111000001011110    0111000001011111    0111000001100000    0111000001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28765 - 28769

  --0111000001100010    0111000001100011    0111000001100100    0111000001100101    0111000001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28770 - 28774

  --0111000001100111    0111000001101000    0111000001101001    0111000001101010    0111000001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28775 - 28779

  --0111000001101100    0111000001101101    0111000001101110    0111000001101111    0111000001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28780 - 28784

  --0111000001110001    0111000001110010    0111000001110011    0111000001110100    0111000001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28785 - 28789

  --0111000001110110    0111000001110111    0111000001111000    0111000001111001    0111000001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28790 - 28794

  --0111000001111011    0111000001111100    0111000001111101    0111000001111110    0111000001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28795 - 28799

  --0111000010000000    0111000010000001    0111000010000010    0111000010000011    0111000010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28800 - 28804

  --0111000010000101    0111000010000110    0111000010000111    0111000010001000    0111000010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28805 - 28809

  --0111000010001010    0111000010001011    0111000010001100    0111000010001101    0111000010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28810 - 28814

  --0111000010001111    0111000010010000    0111000010010001    0111000010010010    0111000010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28815 - 28819

  --0111000010010100    0111000010010101    0111000010010110    0111000010010111    0111000010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28820 - 28824

  --0111000010011001    0111000010011010    0111000010011011    0111000010011100    0111000010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28825 - 28829

  --0111000010011110    0111000010011111    0111000010100000    0111000010100001    0111000010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28830 - 28834

  --0111000010100011    0111000010100100    0111000010100101    0111000010100110    0111000010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28835 - 28839

  --0111000010101000    0111000010101001    0111000010101010    0111000010101011    0111000010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28840 - 28844

  --0111000010101101    0111000010101110    0111000010101111    0111000010110000    0111000010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28845 - 28849

  --0111000010110010    0111000010110011    0111000010110100    0111000010110101    0111000010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28850 - 28854

  --0111000010110111    0111000010111000    0111000010111001    0111000010111010    0111000010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28855 - 28859

  --0111000010111100    0111000010111101    0111000010111110    0111000010111111    0111000011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28860 - 28864

  --0111000011000001    0111000011000010    0111000011000011    0111000011000100    0111000011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28865 - 28869

  --0111000011000110    0111000011000111    0111000011001000    0111000011001001    0111000011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28870 - 28874

  --0111000011001011    0111000011001100    0111000011001101    0111000011001110    0111000011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28875 - 28879

  --0111000011010000    0111000011010001    0111000011010010    0111000011010011    0111000011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28880 - 28884

  --0111000011010101    0111000011010110    0111000011010111    0111000011011000    0111000011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28885 - 28889

  --0111000011011010    0111000011011011    0111000011011100    0111000011011101    0111000011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28890 - 28894

  --0111000011011111    0111000011100000    0111000011100001    0111000011100010    0111000011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28895 - 28899

  --0111000011100100    0111000011100101    0111000011100110    0111000011100111    0111000011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28900 - 28904

  --0111000011101001    0111000011101010    0111000011101011    0111000011101100    0111000011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28905 - 28909

  --0111000011101110    0111000011101111    0111000011110000    0111000011110001    0111000011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28910 - 28914

  --0111000011110011    0111000011110100    0111000011110101    0111000011110110    0111000011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28915 - 28919

  --0111000011111000    0111000011111001    0111000011111010    0111000011111011    0111000011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28920 - 28924

  --0111000011111101    0111000011111110    0111000011111111    0111000100000000    0111000100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28925 - 28929

  --0111000100000010    0111000100000011    0111000100000100    0111000100000101    0111000100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28930 - 28934

  --0111000100000111    0111000100001000    0111000100001001    0111000100001010    0111000100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28935 - 28939

  --0111000100001100    0111000100001101    0111000100001110    0111000100001111    0111000100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28940 - 28944

  --0111000100010001    0111000100010010    0111000100010011    0111000100010100    0111000100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28945 - 28949

  --0111000100010110    0111000100010111    0111000100011000    0111000100011001    0111000100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28950 - 28954

  --0111000100011011    0111000100011100    0111000100011101    0111000100011110    0111000100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28955 - 28959

  --0111000100100000    0111000100100001    0111000100100010    0111000100100011    0111000100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28960 - 28964

  --0111000100100101    0111000100100110    0111000100100111    0111000100101000    0111000100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28965 - 28969

  --0111000100101010    0111000100101011    0111000100101100    0111000100101101    0111000100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28970 - 28974

  --0111000100101111    0111000100110000    0111000100110001    0111000100110010    0111000100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28975 - 28979

  --0111000100110100    0111000100110101    0111000100110110    0111000100110111    0111000100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28980 - 28984

  --0111000100111001    0111000100111010    0111000100111011    0111000100111100    0111000100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28985 - 28989

  --0111000100111110    0111000100111111    0111000101000000    0111000101000001    0111000101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28990 - 28994

  --0111000101000011    0111000101000100    0111000101000101    0111000101000110    0111000101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 28995 - 28999

  --0111000101001000    0111000101001001    0111000101001010    0111000101001011    0111000101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29000 - 29004

  --0111000101001101    0111000101001110    0111000101001111    0111000101010000    0111000101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29005 - 29009

  --0111000101010010    0111000101010011    0111000101010100    0111000101010101    0111000101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29010 - 29014

  --0111000101010111    0111000101011000    0111000101011001    0111000101011010    0111000101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29015 - 29019

  --0111000101011100    0111000101011101    0111000101011110    0111000101011111    0111000101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29020 - 29024

  --0111000101100001    0111000101100010    0111000101100011    0111000101100100    0111000101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29025 - 29029

  --0111000101100110    0111000101100111    0111000101101000    0111000101101001    0111000101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29030 - 29034

  --0111000101101011    0111000101101100    0111000101101101    0111000101101110    0111000101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29035 - 29039

  --0111000101110000    0111000101110001    0111000101110010    0111000101110011    0111000101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29040 - 29044

  --0111000101110101    0111000101110110    0111000101110111    0111000101111000    0111000101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29045 - 29049

  --0111000101111010    0111000101111011    0111000101111100    0111000101111101    0111000101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29050 - 29054

  --0111000101111111    0111000110000000    0111000110000001    0111000110000010    0111000110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29055 - 29059

  --0111000110000100    0111000110000101    0111000110000110    0111000110000111    0111000110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29060 - 29064

  --0111000110001001    0111000110001010    0111000110001011    0111000110001100    0111000110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29065 - 29069

  --0111000110001110    0111000110001111    0111000110010000    0111000110010001    0111000110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29070 - 29074

  --0111000110010011    0111000110010100    0111000110010101    0111000110010110    0111000110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29075 - 29079

  --0111000110011000    0111000110011001    0111000110011010    0111000110011011    0111000110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29080 - 29084

  --0111000110011101    0111000110011110    0111000110011111    0111000110100000    0111000110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29085 - 29089

  --0111000110100010    0111000110100011    0111000110100100    0111000110100101    0111000110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29090 - 29094

  --0111000110100111    0111000110101000    0111000110101001    0111000110101010    0111000110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29095 - 29099

  --0111000110101100    0111000110101101    0111000110101110    0111000110101111    0111000110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29100 - 29104

  --0111000110110001    0111000110110010    0111000110110011    0111000110110100    0111000110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29105 - 29109

  --0111000110110110    0111000110110111    0111000110111000    0111000110111001    0111000110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29110 - 29114

  --0111000110111011    0111000110111100    0111000110111101    0111000110111110    0111000110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29115 - 29119

  --0111000111000000    0111000111000001    0111000111000010    0111000111000011    0111000111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29120 - 29124

  --0111000111000101    0111000111000110    0111000111000111    0111000111001000    0111000111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29125 - 29129

  --0111000111001010    0111000111001011    0111000111001100    0111000111001101    0111000111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29130 - 29134

  --0111000111001111    0111000111010000    0111000111010001    0111000111010010    0111000111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29135 - 29139

  --0111000111010100    0111000111010101    0111000111010110    0111000111010111    0111000111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29140 - 29144

  --0111000111011001    0111000111011010    0111000111011011    0111000111011100    0111000111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29145 - 29149

  --0111000111011110    0111000111011111    0111000111100000    0111000111100001    0111000111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29150 - 29154

  --0111000111100011    0111000111100100    0111000111100101    0111000111100110    0111000111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29155 - 29159

  --0111000111101000    0111000111101001    0111000111101010    0111000111101011    0111000111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29160 - 29164

  --0111000111101101    0111000111101110    0111000111101111    0111000111110000    0111000111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29165 - 29169

  --0111000111110010    0111000111110011    0111000111110100    0111000111110101    0111000111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29170 - 29174

  --0111000111110111    0111000111111000    0111000111111001    0111000111111010    0111000111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29175 - 29179

  --0111000111111100    0111000111111101    0111000111111110    0111000111111111    0111001000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29180 - 29184

  --0111001000000001    0111001000000010    0111001000000011    0111001000000100    0111001000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29185 - 29189

  --0111001000000110    0111001000000111    0111001000001000    0111001000001001    0111001000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29190 - 29194

  --0111001000001011    0111001000001100    0111001000001101    0111001000001110    0111001000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29195 - 29199

  --0111001000010000    0111001000010001    0111001000010010    0111001000010011    0111001000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29200 - 29204

  --0111001000010101    0111001000010110    0111001000010111    0111001000011000    0111001000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29205 - 29209

  --0111001000011010    0111001000011011    0111001000011100    0111001000011101    0111001000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29210 - 29214

  --0111001000011111    0111001000100000    0111001000100001    0111001000100010    0111001000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29215 - 29219

  --0111001000100100    0111001000100101    0111001000100110    0111001000100111    0111001000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29220 - 29224

  --0111001000101001    0111001000101010    0111001000101011    0111001000101100    0111001000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29225 - 29229

  --0111001000101110    0111001000101111    0111001000110000    0111001000110001    0111001000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29230 - 29234

  --0111001000110011    0111001000110100    0111001000110101    0111001000110110    0111001000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29235 - 29239

  --0111001000111000    0111001000111001    0111001000111010    0111001000111011    0111001000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29240 - 29244

  --0111001000111101    0111001000111110    0111001000111111    0111001001000000    0111001001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29245 - 29249

  --0111001001000010    0111001001000011    0111001001000100    0111001001000101    0111001001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29250 - 29254

  --0111001001000111    0111001001001000    0111001001001001    0111001001001010    0111001001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29255 - 29259

  --0111001001001100    0111001001001101    0111001001001110    0111001001001111    0111001001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29260 - 29264

  --0111001001010001    0111001001010010    0111001001010011    0111001001010100    0111001001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29265 - 29269

  --0111001001010110    0111001001010111    0111001001011000    0111001001011001    0111001001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29270 - 29274

  --0111001001011011    0111001001011100    0111001001011101    0111001001011110    0111001001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29275 - 29279

  --0111001001100000    0111001001100001    0111001001100010    0111001001100011    0111001001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29280 - 29284

  --0111001001100101    0111001001100110    0111001001100111    0111001001101000    0111001001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29285 - 29289

  --0111001001101010    0111001001101011    0111001001101100    0111001001101101    0111001001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29290 - 29294

  --0111001001101111    0111001001110000    0111001001110001    0111001001110010    0111001001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29295 - 29299

  --0111001001110100    0111001001110101    0111001001110110    0111001001110111    0111001001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29300 - 29304

  --0111001001111001    0111001001111010    0111001001111011    0111001001111100    0111001001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29305 - 29309

  --0111001001111110    0111001001111111    0111001010000000    0111001010000001    0111001010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29310 - 29314

  --0111001010000011    0111001010000100    0111001010000101    0111001010000110    0111001010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29315 - 29319

  --0111001010001000    0111001010001001    0111001010001010    0111001010001011    0111001010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29320 - 29324

  --0111001010001101    0111001010001110    0111001010001111    0111001010010000    0111001010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29325 - 29329

  --0111001010010010    0111001010010011    0111001010010100    0111001010010101    0111001010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29330 - 29334

  --0111001010010111    0111001010011000    0111001010011001    0111001010011010    0111001010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29335 - 29339

  --0111001010011100    0111001010011101    0111001010011110    0111001010011111    0111001010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29340 - 29344

  --0111001010100001    0111001010100010    0111001010100011    0111001010100100    0111001010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29345 - 29349

  --0111001010100110    0111001010100111    0111001010101000    0111001010101001    0111001010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29350 - 29354

  --0111001010101011    0111001010101100    0111001010101101    0111001010101110    0111001010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29355 - 29359

  --0111001010110000    0111001010110001    0111001010110010    0111001010110011    0111001010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29360 - 29364

  --0111001010110101    0111001010110110    0111001010110111    0111001010111000    0111001010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29365 - 29369

  --0111001010111010    0111001010111011    0111001010111100    0111001010111101    0111001010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29370 - 29374

  --0111001010111111    0111001011000000    0111001011000001    0111001011000010    0111001011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29375 - 29379

  --0111001011000100    0111001011000101    0111001011000110    0111001011000111    0111001011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29380 - 29384

  --0111001011001001    0111001011001010    0111001011001011    0111001011001100    0111001011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29385 - 29389

  --0111001011001110    0111001011001111    0111001011010000    0111001011010001    0111001011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29390 - 29394

  --0111001011010011    0111001011010100    0111001011010101    0111001011010110    0111001011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29395 - 29399

  --0111001011011000    0111001011011001    0111001011011010    0111001011011011    0111001011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29400 - 29404

  --0111001011011101    0111001011011110    0111001011011111    0111001011100000    0111001011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29405 - 29409

  --0111001011100010    0111001011100011    0111001011100100    0111001011100101    0111001011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29410 - 29414

  --0111001011100111    0111001011101000    0111001011101001    0111001011101010    0111001011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29415 - 29419

  --0111001011101100    0111001011101101    0111001011101110    0111001011101111    0111001011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29420 - 29424

  --0111001011110001    0111001011110010    0111001011110011    0111001011110100    0111001011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29425 - 29429

  --0111001011110110    0111001011110111    0111001011111000    0111001011111001    0111001011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29430 - 29434

  --0111001011111011    0111001011111100    0111001011111101    0111001011111110    0111001011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29435 - 29439

  --0111001100000000    0111001100000001    0111001100000010    0111001100000011    0111001100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29440 - 29444

  --0111001100000101    0111001100000110    0111001100000111    0111001100001000    0111001100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29445 - 29449

  --0111001100001010    0111001100001011    0111001100001100    0111001100001101    0111001100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29450 - 29454

  --0111001100001111    0111001100010000    0111001100010001    0111001100010010    0111001100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29455 - 29459

  --0111001100010100    0111001100010101    0111001100010110    0111001100010111    0111001100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29460 - 29464

  --0111001100011001    0111001100011010    0111001100011011    0111001100011100    0111001100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29465 - 29469

  --0111001100011110    0111001100011111    0111001100100000    0111001100100001    0111001100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29470 - 29474

  --0111001100100011    0111001100100100    0111001100100101    0111001100100110    0111001100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29475 - 29479

  --0111001100101000    0111001100101001    0111001100101010    0111001100101011    0111001100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29480 - 29484

  --0111001100101101    0111001100101110    0111001100101111    0111001100110000    0111001100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29485 - 29489

  --0111001100110010    0111001100110011    0111001100110100    0111001100110101    0111001100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29490 - 29494

  --0111001100110111    0111001100111000    0111001100111001    0111001100111010    0111001100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29495 - 29499

  --0111001100111100    0111001100111101    0111001100111110    0111001100111111    0111001101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29500 - 29504

  --0111001101000001    0111001101000010    0111001101000011    0111001101000100    0111001101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29505 - 29509

  --0111001101000110    0111001101000111    0111001101001000    0111001101001001    0111001101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29510 - 29514

  --0111001101001011    0111001101001100    0111001101001101    0111001101001110    0111001101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29515 - 29519

  --0111001101010000    0111001101010001    0111001101010010    0111001101010011    0111001101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29520 - 29524

  --0111001101010101    0111001101010110    0111001101010111    0111001101011000    0111001101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29525 - 29529

  --0111001101011010    0111001101011011    0111001101011100    0111001101011101    0111001101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29530 - 29534

  --0111001101011111    0111001101100000    0111001101100001    0111001101100010    0111001101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29535 - 29539

  --0111001101100100    0111001101100101    0111001101100110    0111001101100111    0111001101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29540 - 29544

  --0111001101101001    0111001101101010    0111001101101011    0111001101101100    0111001101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29545 - 29549

  --0111001101101110    0111001101101111    0111001101110000    0111001101110001    0111001101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29550 - 29554

  --0111001101110011    0111001101110100    0111001101110101    0111001101110110    0111001101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29555 - 29559

  --0111001101111000    0111001101111001    0111001101111010    0111001101111011    0111001101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29560 - 29564

  --0111001101111101    0111001101111110    0111001101111111    0111001110000000    0111001110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29565 - 29569

  --0111001110000010    0111001110000011    0111001110000100    0111001110000101    0111001110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29570 - 29574

  --0111001110000111    0111001110001000    0111001110001001    0111001110001010    0111001110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29575 - 29579

  --0111001110001100    0111001110001101    0111001110001110    0111001110001111    0111001110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29580 - 29584

  --0111001110010001    0111001110010010    0111001110010011    0111001110010100    0111001110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29585 - 29589

  --0111001110010110    0111001110010111    0111001110011000    0111001110011001    0111001110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29590 - 29594

  --0111001110011011    0111001110011100    0111001110011101    0111001110011110    0111001110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29595 - 29599

  --0111001110100000    0111001110100001    0111001110100010    0111001110100011    0111001110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29600 - 29604

  --0111001110100101    0111001110100110    0111001110100111    0111001110101000    0111001110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29605 - 29609

  --0111001110101010    0111001110101011    0111001110101100    0111001110101101    0111001110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29610 - 29614

  --0111001110101111    0111001110110000    0111001110110001    0111001110110010    0111001110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29615 - 29619

  --0111001110110100    0111001110110101    0111001110110110    0111001110110111    0111001110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29620 - 29624

  --0111001110111001    0111001110111010    0111001110111011    0111001110111100    0111001110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29625 - 29629

  --0111001110111110    0111001110111111    0111001111000000    0111001111000001    0111001111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29630 - 29634

  --0111001111000011    0111001111000100    0111001111000101    0111001111000110    0111001111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29635 - 29639

  --0111001111001000    0111001111001001    0111001111001010    0111001111001011    0111001111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29640 - 29644

  --0111001111001101    0111001111001110    0111001111001111    0111001111010000    0111001111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29645 - 29649

  --0111001111010010    0111001111010011    0111001111010100    0111001111010101    0111001111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29650 - 29654

  --0111001111010111    0111001111011000    0111001111011001    0111001111011010    0111001111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29655 - 29659

  --0111001111011100    0111001111011101    0111001111011110    0111001111011111    0111001111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29660 - 29664

  --0111001111100001    0111001111100010    0111001111100011    0111001111100100    0111001111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29665 - 29669

  --0111001111100110    0111001111100111    0111001111101000    0111001111101001    0111001111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29670 - 29674

  --0111001111101011    0111001111101100    0111001111101101    0111001111101110    0111001111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29675 - 29679

  --0111001111110000    0111001111110001    0111001111110010    0111001111110011    0111001111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29680 - 29684

  --0111001111110101    0111001111110110    0111001111110111    0111001111111000    0111001111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29685 - 29689

  --0111001111111010    0111001111111011    0111001111111100    0111001111111101    0111001111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29690 - 29694

  --0111001111111111    0111010000000000    0111010000000001    0111010000000010    0111010000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29695 - 29699

  --0111010000000100    0111010000000101    0111010000000110    0111010000000111    0111010000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29700 - 29704

  --0111010000001001    0111010000001010    0111010000001011    0111010000001100    0111010000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29705 - 29709

  --0111010000001110    0111010000001111    0111010000010000    0111010000010001    0111010000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29710 - 29714

  --0111010000010011    0111010000010100    0111010000010101    0111010000010110    0111010000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29715 - 29719

  --0111010000011000    0111010000011001    0111010000011010    0111010000011011    0111010000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29720 - 29724

  --0111010000011101    0111010000011110    0111010000011111    0111010000100000    0111010000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29725 - 29729

  --0111010000100010    0111010000100011    0111010000100100    0111010000100101    0111010000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29730 - 29734

  --0111010000100111    0111010000101000    0111010000101001    0111010000101010    0111010000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29735 - 29739

  --0111010000101100    0111010000101101    0111010000101110    0111010000101111    0111010000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29740 - 29744

  --0111010000110001    0111010000110010    0111010000110011    0111010000110100    0111010000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29745 - 29749

  --0111010000110110    0111010000110111    0111010000111000    0111010000111001    0111010000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29750 - 29754

  --0111010000111011    0111010000111100    0111010000111101    0111010000111110    0111010000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29755 - 29759

  --0111010001000000    0111010001000001    0111010001000010    0111010001000011    0111010001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29760 - 29764

  --0111010001000101    0111010001000110    0111010001000111    0111010001001000    0111010001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29765 - 29769

  --0111010001001010    0111010001001011    0111010001001100    0111010001001101    0111010001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29770 - 29774

  --0111010001001111    0111010001010000    0111010001010001    0111010001010010    0111010001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29775 - 29779

  --0111010001010100    0111010001010101    0111010001010110    0111010001010111    0111010001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29780 - 29784

  --0111010001011001    0111010001011010    0111010001011011    0111010001011100    0111010001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29785 - 29789

  --0111010001011110    0111010001011111    0111010001100000    0111010001100001    0111010001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29790 - 29794

  --0111010001100011    0111010001100100    0111010001100101    0111010001100110    0111010001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29795 - 29799

  --0111010001101000    0111010001101001    0111010001101010    0111010001101011    0111010001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29800 - 29804

  --0111010001101101    0111010001101110    0111010001101111    0111010001110000    0111010001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29805 - 29809

  --0111010001110010    0111010001110011    0111010001110100    0111010001110101    0111010001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29810 - 29814

  --0111010001110111    0111010001111000    0111010001111001    0111010001111010    0111010001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29815 - 29819

  --0111010001111100    0111010001111101    0111010001111110    0111010001111111    0111010010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29820 - 29824

  --0111010010000001    0111010010000010    0111010010000011    0111010010000100    0111010010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29825 - 29829

  --0111010010000110    0111010010000111    0111010010001000    0111010010001001    0111010010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29830 - 29834

  --0111010010001011    0111010010001100    0111010010001101    0111010010001110    0111010010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29835 - 29839

  --0111010010010000    0111010010010001    0111010010010010    0111010010010011    0111010010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29840 - 29844

  --0111010010010101    0111010010010110    0111010010010111    0111010010011000    0111010010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29845 - 29849

  --0111010010011010    0111010010011011    0111010010011100    0111010010011101    0111010010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29850 - 29854

  --0111010010011111    0111010010100000    0111010010100001    0111010010100010    0111010010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29855 - 29859

  --0111010010100100    0111010010100101    0111010010100110    0111010010100111    0111010010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29860 - 29864

  --0111010010101001    0111010010101010    0111010010101011    0111010010101100    0111010010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29865 - 29869

  --0111010010101110    0111010010101111    0111010010110000    0111010010110001    0111010010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29870 - 29874

  --0111010010110011    0111010010110100    0111010010110101    0111010010110110    0111010010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29875 - 29879

  --0111010010111000    0111010010111001    0111010010111010    0111010010111011    0111010010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29880 - 29884

  --0111010010111101    0111010010111110    0111010010111111    0111010011000000    0111010011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29885 - 29889

  --0111010011000010    0111010011000011    0111010011000100    0111010011000101    0111010011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29890 - 29894

  --0111010011000111    0111010011001000    0111010011001001    0111010011001010    0111010011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29895 - 29899

  --0111010011001100    0111010011001101    0111010011001110    0111010011001111    0111010011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29900 - 29904

  --0111010011010001    0111010011010010    0111010011010011    0111010011010100    0111010011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29905 - 29909

  --0111010011010110    0111010011010111    0111010011011000    0111010011011001    0111010011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29910 - 29914

  --0111010011011011    0111010011011100    0111010011011101    0111010011011110    0111010011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29915 - 29919

  --0111010011100000    0111010011100001    0111010011100010    0111010011100011    0111010011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29920 - 29924

  --0111010011100101    0111010011100110    0111010011100111    0111010011101000    0111010011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29925 - 29929

  --0111010011101010    0111010011101011    0111010011101100    0111010011101101    0111010011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29930 - 29934

  --0111010011101111    0111010011110000    0111010011110001    0111010011110010    0111010011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29935 - 29939

  --0111010011110100    0111010011110101    0111010011110110    0111010011110111    0111010011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29940 - 29944

  --0111010011111001    0111010011111010    0111010011111011    0111010011111100    0111010011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29945 - 29949

  --0111010011111110    0111010011111111    0111010100000000    0111010100000001    0111010100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29950 - 29954

  --0111010100000011    0111010100000100    0111010100000101    0111010100000110    0111010100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29955 - 29959

  --0111010100001000    0111010100001001    0111010100001010    0111010100001011    0111010100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29960 - 29964

  --0111010100001101    0111010100001110    0111010100001111    0111010100010000    0111010100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29965 - 29969

  --0111010100010010    0111010100010011    0111010100010100    0111010100010101    0111010100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29970 - 29974

  --0111010100010111    0111010100011000    0111010100011001    0111010100011010    0111010100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29975 - 29979

  --0111010100011100    0111010100011101    0111010100011110    0111010100011111    0111010100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29980 - 29984

  --0111010100100001    0111010100100010    0111010100100011    0111010100100100    0111010100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29985 - 29989

  --0111010100100110    0111010100100111    0111010100101000    0111010100101001    0111010100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29990 - 29994

  --0111010100101011    0111010100101100    0111010100101101    0111010100101110    0111010100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 29995 - 29999

  --0111010100110000    0111010100110001    0111010100110010    0111010100110011    0111010100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30000 - 30004

  --0111010100110101    0111010100110110    0111010100110111    0111010100111000    0111010100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30005 - 30009

  --0111010100111010    0111010100111011    0111010100111100    0111010100111101    0111010100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30010 - 30014

  --0111010100111111    0111010101000000    0111010101000001    0111010101000010    0111010101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30015 - 30019

  --0111010101000100    0111010101000101    0111010101000110    0111010101000111    0111010101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30020 - 30024

  --0111010101001001    0111010101001010    0111010101001011    0111010101001100    0111010101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30025 - 30029

  --0111010101001110    0111010101001111    0111010101010000    0111010101010001    0111010101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30030 - 30034

  --0111010101010011    0111010101010100    0111010101010101    0111010101010110    0111010101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30035 - 30039

  --0111010101011000    0111010101011001    0111010101011010    0111010101011011    0111010101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30040 - 30044

  --0111010101011101    0111010101011110    0111010101011111    0111010101100000    0111010101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30045 - 30049

  --0111010101100010    0111010101100011    0111010101100100    0111010101100101    0111010101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30050 - 30054

  --0111010101100111    0111010101101000    0111010101101001    0111010101101010    0111010101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30055 - 30059

  --0111010101101100    0111010101101101    0111010101101110    0111010101101111    0111010101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30060 - 30064

  --0111010101110001    0111010101110010    0111010101110011    0111010101110100    0111010101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30065 - 30069

  --0111010101110110    0111010101110111    0111010101111000    0111010101111001    0111010101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30070 - 30074

  --0111010101111011    0111010101111100    0111010101111101    0111010101111110    0111010101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30075 - 30079

  --0111010110000000    0111010110000001    0111010110000010    0111010110000011    0111010110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30080 - 30084

  --0111010110000101    0111010110000110    0111010110000111    0111010110001000    0111010110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30085 - 30089

  --0111010110001010    0111010110001011    0111010110001100    0111010110001101    0111010110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30090 - 30094

  --0111010110001111    0111010110010000    0111010110010001    0111010110010010    0111010110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30095 - 30099

  --0111010110010100    0111010110010101    0111010110010110    0111010110010111    0111010110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30100 - 30104

  --0111010110011001    0111010110011010    0111010110011011    0111010110011100    0111010110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30105 - 30109

  --0111010110011110    0111010110011111    0111010110100000    0111010110100001    0111010110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30110 - 30114

  --0111010110100011    0111010110100100    0111010110100101    0111010110100110    0111010110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30115 - 30119

  --0111010110101000    0111010110101001    0111010110101010    0111010110101011    0111010110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30120 - 30124

  --0111010110101101    0111010110101110    0111010110101111    0111010110110000    0111010110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30125 - 30129

  --0111010110110010    0111010110110011    0111010110110100    0111010110110101    0111010110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30130 - 30134

  --0111010110110111    0111010110111000    0111010110111001    0111010110111010    0111010110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30135 - 30139

  --0111010110111100    0111010110111101    0111010110111110    0111010110111111    0111010111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30140 - 30144

  --0111010111000001    0111010111000010    0111010111000011    0111010111000100    0111010111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30145 - 30149

  --0111010111000110    0111010111000111    0111010111001000    0111010111001001    0111010111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30150 - 30154

  --0111010111001011    0111010111001100    0111010111001101    0111010111001110    0111010111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30155 - 30159

  --0111010111010000    0111010111010001    0111010111010010    0111010111010011    0111010111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30160 - 30164

  --0111010111010101    0111010111010110    0111010111010111    0111010111011000    0111010111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30165 - 30169

  --0111010111011010    0111010111011011    0111010111011100    0111010111011101    0111010111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30170 - 30174

  --0111010111011111    0111010111100000    0111010111100001    0111010111100010    0111010111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30175 - 30179

  --0111010111100100    0111010111100101    0111010111100110    0111010111100111    0111010111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30180 - 30184

  --0111010111101001    0111010111101010    0111010111101011    0111010111101100    0111010111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30185 - 30189

  --0111010111101110    0111010111101111    0111010111110000    0111010111110001    0111010111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30190 - 30194

  --0111010111110011    0111010111110100    0111010111110101    0111010111110110    0111010111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30195 - 30199

  --0111010111111000    0111010111111001    0111010111111010    0111010111111011    0111010111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30200 - 30204

  --0111010111111101    0111010111111110    0111010111111111    0111011000000000    0111011000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30205 - 30209

  --0111011000000010    0111011000000011    0111011000000100    0111011000000101    0111011000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30210 - 30214

  --0111011000000111    0111011000001000    0111011000001001    0111011000001010    0111011000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30215 - 30219

  --0111011000001100    0111011000001101    0111011000001110    0111011000001111    0111011000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30220 - 30224

  --0111011000010001    0111011000010010    0111011000010011    0111011000010100    0111011000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30225 - 30229

  --0111011000010110    0111011000010111    0111011000011000    0111011000011001    0111011000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30230 - 30234

  --0111011000011011    0111011000011100    0111011000011101    0111011000011110    0111011000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30235 - 30239

  --0111011000100000    0111011000100001    0111011000100010    0111011000100011    0111011000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30240 - 30244

  --0111011000100101    0111011000100110    0111011000100111    0111011000101000    0111011000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30245 - 30249

  --0111011000101010    0111011000101011    0111011000101100    0111011000101101    0111011000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30250 - 30254

  --0111011000101111    0111011000110000    0111011000110001    0111011000110010    0111011000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30255 - 30259

  --0111011000110100    0111011000110101    0111011000110110    0111011000110111    0111011000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30260 - 30264

  --0111011000111001    0111011000111010    0111011000111011    0111011000111100    0111011000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30265 - 30269

  --0111011000111110    0111011000111111    0111011001000000    0111011001000001    0111011001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30270 - 30274

  --0111011001000011    0111011001000100    0111011001000101    0111011001000110    0111011001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30275 - 30279

  --0111011001001000    0111011001001001    0111011001001010    0111011001001011    0111011001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30280 - 30284

  --0111011001001101    0111011001001110    0111011001001111    0111011001010000    0111011001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30285 - 30289

  --0111011001010010    0111011001010011    0111011001010100    0111011001010101    0111011001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30290 - 30294

  --0111011001010111    0111011001011000    0111011001011001    0111011001011010    0111011001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30295 - 30299

  --0111011001011100    0111011001011101    0111011001011110    0111011001011111    0111011001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30300 - 30304

  --0111011001100001    0111011001100010    0111011001100011    0111011001100100    0111011001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30305 - 30309

  --0111011001100110    0111011001100111    0111011001101000    0111011001101001    0111011001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30310 - 30314

  --0111011001101011    0111011001101100    0111011001101101    0111011001101110    0111011001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30315 - 30319

  --0111011001110000    0111011001110001    0111011001110010    0111011001110011    0111011001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30320 - 30324

  --0111011001110101    0111011001110110    0111011001110111    0111011001111000    0111011001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30325 - 30329

  --0111011001111010    0111011001111011    0111011001111100    0111011001111101    0111011001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30330 - 30334

  --0111011001111111    0111011010000000    0111011010000001    0111011010000010    0111011010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30335 - 30339

  --0111011010000100    0111011010000101    0111011010000110    0111011010000111    0111011010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30340 - 30344

  --0111011010001001    0111011010001010    0111011010001011    0111011010001100    0111011010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30345 - 30349

  --0111011010001110    0111011010001111    0111011010010000    0111011010010001    0111011010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30350 - 30354

  --0111011010010011    0111011010010100    0111011010010101    0111011010010110    0111011010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30355 - 30359

  --0111011010011000    0111011010011001    0111011010011010    0111011010011011    0111011010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30360 - 30364

  --0111011010011101    0111011010011110    0111011010011111    0111011010100000    0111011010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30365 - 30369

  --0111011010100010    0111011010100011    0111011010100100    0111011010100101    0111011010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30370 - 30374

  --0111011010100111    0111011010101000    0111011010101001    0111011010101010    0111011010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30375 - 30379

  --0111011010101100    0111011010101101    0111011010101110    0111011010101111    0111011010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30380 - 30384

  --0111011010110001    0111011010110010    0111011010110011    0111011010110100    0111011010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30385 - 30389

  --0111011010110110    0111011010110111    0111011010111000    0111011010111001    0111011010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30390 - 30394

  --0111011010111011    0111011010111100    0111011010111101    0111011010111110    0111011010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30395 - 30399

  --0111011011000000    0111011011000001    0111011011000010    0111011011000011    0111011011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30400 - 30404

  --0111011011000101    0111011011000110    0111011011000111    0111011011001000    0111011011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30405 - 30409

  --0111011011001010    0111011011001011    0111011011001100    0111011011001101    0111011011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30410 - 30414

  --0111011011001111    0111011011010000    0111011011010001    0111011011010010    0111011011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30415 - 30419

  --0111011011010100    0111011011010101    0111011011010110    0111011011010111    0111011011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30420 - 30424

  --0111011011011001    0111011011011010    0111011011011011    0111011011011100    0111011011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30425 - 30429

  --0111011011011110    0111011011011111    0111011011100000    0111011011100001    0111011011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30430 - 30434

  --0111011011100011    0111011011100100    0111011011100101    0111011011100110    0111011011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30435 - 30439

  --0111011011101000    0111011011101001    0111011011101010    0111011011101011    0111011011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30440 - 30444

  --0111011011101101    0111011011101110    0111011011101111    0111011011110000    0111011011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30445 - 30449

  --0111011011110010    0111011011110011    0111011011110100    0111011011110101    0111011011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30450 - 30454

  --0111011011110111    0111011011111000    0111011011111001    0111011011111010    0111011011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30455 - 30459

  --0111011011111100    0111011011111101    0111011011111110    0111011011111111    0111011100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30460 - 30464

  --0111011100000001    0111011100000010    0111011100000011    0111011100000100    0111011100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30465 - 30469

  --0111011100000110    0111011100000111    0111011100001000    0111011100001001    0111011100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30470 - 30474

  --0111011100001011    0111011100001100    0111011100001101    0111011100001110    0111011100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30475 - 30479

  --0111011100010000    0111011100010001    0111011100010010    0111011100010011    0111011100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30480 - 30484

  --0111011100010101    0111011100010110    0111011100010111    0111011100011000    0111011100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30485 - 30489

  --0111011100011010    0111011100011011    0111011100011100    0111011100011101    0111011100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30490 - 30494

  --0111011100011111    0111011100100000    0111011100100001    0111011100100010    0111011100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30495 - 30499

  --0111011100100100    0111011100100101    0111011100100110    0111011100100111    0111011100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30500 - 30504

  --0111011100101001    0111011100101010    0111011100101011    0111011100101100    0111011100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30505 - 30509

  --0111011100101110    0111011100101111    0111011100110000    0111011100110001    0111011100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30510 - 30514

  --0111011100110011    0111011100110100    0111011100110101    0111011100110110    0111011100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30515 - 30519

  --0111011100111000    0111011100111001    0111011100111010    0111011100111011    0111011100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30520 - 30524

  --0111011100111101    0111011100111110    0111011100111111    0111011101000000    0111011101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30525 - 30529

  --0111011101000010    0111011101000011    0111011101000100    0111011101000101    0111011101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30530 - 30534

  --0111011101000111    0111011101001000    0111011101001001    0111011101001010    0111011101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30535 - 30539

  --0111011101001100    0111011101001101    0111011101001110    0111011101001111    0111011101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30540 - 30544

  --0111011101010001    0111011101010010    0111011101010011    0111011101010100    0111011101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30545 - 30549

  --0111011101010110    0111011101010111    0111011101011000    0111011101011001    0111011101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30550 - 30554

  --0111011101011011    0111011101011100    0111011101011101    0111011101011110    0111011101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30555 - 30559

  --0111011101100000    0111011101100001    0111011101100010    0111011101100011    0111011101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30560 - 30564

  --0111011101100101    0111011101100110    0111011101100111    0111011101101000    0111011101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30565 - 30569

  --0111011101101010    0111011101101011    0111011101101100    0111011101101101    0111011101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30570 - 30574

  --0111011101101111    0111011101110000    0111011101110001    0111011101110010    0111011101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30575 - 30579

  --0111011101110100    0111011101110101    0111011101110110    0111011101110111    0111011101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30580 - 30584

  --0111011101111001    0111011101111010    0111011101111011    0111011101111100    0111011101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30585 - 30589

  --0111011101111110    0111011101111111    0111011110000000    0111011110000001    0111011110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30590 - 30594

  --0111011110000011    0111011110000100    0111011110000101    0111011110000110    0111011110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30595 - 30599

  --0111011110001000    0111011110001001    0111011110001010    0111011110001011    0111011110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30600 - 30604

  --0111011110001101    0111011110001110    0111011110001111    0111011110010000    0111011110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30605 - 30609

  --0111011110010010    0111011110010011    0111011110010100    0111011110010101    0111011110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30610 - 30614

  --0111011110010111    0111011110011000    0111011110011001    0111011110011010    0111011110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30615 - 30619

  --0111011110011100    0111011110011101    0111011110011110    0111011110011111    0111011110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30620 - 30624

  --0111011110100001    0111011110100010    0111011110100011    0111011110100100    0111011110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30625 - 30629

  --0111011110100110    0111011110100111    0111011110101000    0111011110101001    0111011110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30630 - 30634

  --0111011110101011    0111011110101100    0111011110101101    0111011110101110    0111011110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30635 - 30639

  --0111011110110000    0111011110110001    0111011110110010    0111011110110011    0111011110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30640 - 30644

  --0111011110110101    0111011110110110    0111011110110111    0111011110111000    0111011110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30645 - 30649

  --0111011110111010    0111011110111011    0111011110111100    0111011110111101    0111011110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30650 - 30654

  --0111011110111111    0111011111000000    0111011111000001    0111011111000010    0111011111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30655 - 30659

  --0111011111000100    0111011111000101    0111011111000110    0111011111000111    0111011111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30660 - 30664

  --0111011111001001    0111011111001010    0111011111001011    0111011111001100    0111011111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30665 - 30669

  --0111011111001110    0111011111001111    0111011111010000    0111011111010001    0111011111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30670 - 30674

  --0111011111010011    0111011111010100    0111011111010101    0111011111010110    0111011111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30675 - 30679

  --0111011111011000    0111011111011001    0111011111011010    0111011111011011    0111011111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30680 - 30684

  --0111011111011101    0111011111011110    0111011111011111    0111011111100000    0111011111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30685 - 30689

  --0111011111100010    0111011111100011    0111011111100100    0111011111100101    0111011111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30690 - 30694

  --0111011111100111    0111011111101000    0111011111101001    0111011111101010    0111011111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30695 - 30699

  --0111011111101100    0111011111101101    0111011111101110    0111011111101111    0111011111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30700 - 30704

  --0111011111110001    0111011111110010    0111011111110011    0111011111110100    0111011111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30705 - 30709

  --0111011111110110    0111011111110111    0111011111111000    0111011111111001    0111011111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30710 - 30714

  --0111011111111011    0111011111111100    0111011111111101    0111011111111110    0111011111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30715 - 30719

  --0111100000000000    0111100000000001    0111100000000010    0111100000000011    0111100000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30720 - 30724

  --0111100000000101    0111100000000110    0111100000000111    0111100000001000    0111100000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30725 - 30729

  --0111100000001010    0111100000001011    0111100000001100    0111100000001101    0111100000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30730 - 30734

  --0111100000001111    0111100000010000    0111100000010001    0111100000010010    0111100000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30735 - 30739

  --0111100000010100    0111100000010101    0111100000010110    0111100000010111    0111100000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30740 - 30744

  --0111100000011001    0111100000011010    0111100000011011    0111100000011100    0111100000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30745 - 30749

  --0111100000011110    0111100000011111    0111100000100000    0111100000100001    0111100000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30750 - 30754

  --0111100000100011    0111100000100100    0111100000100101    0111100000100110    0111100000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30755 - 30759

  --0111100000101000    0111100000101001    0111100000101010    0111100000101011    0111100000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30760 - 30764

  --0111100000101101    0111100000101110    0111100000101111    0111100000110000    0111100000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30765 - 30769

  --0111100000110010    0111100000110011    0111100000110100    0111100000110101    0111100000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30770 - 30774

  --0111100000110111    0111100000111000    0111100000111001    0111100000111010    0111100000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30775 - 30779

  --0111100000111100    0111100000111101    0111100000111110    0111100000111111    0111100001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30780 - 30784

  --0111100001000001    0111100001000010    0111100001000011    0111100001000100    0111100001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30785 - 30789

  --0111100001000110    0111100001000111    0111100001001000    0111100001001001    0111100001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30790 - 30794

  --0111100001001011    0111100001001100    0111100001001101    0111100001001110    0111100001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30795 - 30799

  --0111100001010000    0111100001010001    0111100001010010    0111100001010011    0111100001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30800 - 30804

  --0111100001010101    0111100001010110    0111100001010111    0111100001011000    0111100001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30805 - 30809

  --0111100001011010    0111100001011011    0111100001011100    0111100001011101    0111100001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30810 - 30814

  --0111100001011111    0111100001100000    0111100001100001    0111100001100010    0111100001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30815 - 30819

  --0111100001100100    0111100001100101    0111100001100110    0111100001100111    0111100001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30820 - 30824

  --0111100001101001    0111100001101010    0111100001101011    0111100001101100    0111100001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30825 - 30829

  --0111100001101110    0111100001101111    0111100001110000    0111100001110001    0111100001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30830 - 30834

  --0111100001110011    0111100001110100    0111100001110101    0111100001110110    0111100001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30835 - 30839

  --0111100001111000    0111100001111001    0111100001111010    0111100001111011    0111100001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30840 - 30844

  --0111100001111101    0111100001111110    0111100001111111    0111100010000000    0111100010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30845 - 30849

  --0111100010000010    0111100010000011    0111100010000100    0111100010000101    0111100010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30850 - 30854

  --0111100010000111    0111100010001000    0111100010001001    0111100010001010    0111100010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30855 - 30859

  --0111100010001100    0111100010001101    0111100010001110    0111100010001111    0111100010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30860 - 30864

  --0111100010010001    0111100010010010    0111100010010011    0111100010010100    0111100010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30865 - 30869

  --0111100010010110    0111100010010111    0111100010011000    0111100010011001    0111100010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30870 - 30874

  --0111100010011011    0111100010011100    0111100010011101    0111100010011110    0111100010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30875 - 30879

  --0111100010100000    0111100010100001    0111100010100010    0111100010100011    0111100010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30880 - 30884

  --0111100010100101    0111100010100110    0111100010100111    0111100010101000    0111100010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30885 - 30889

  --0111100010101010    0111100010101011    0111100010101100    0111100010101101    0111100010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30890 - 30894

  --0111100010101111    0111100010110000    0111100010110001    0111100010110010    0111100010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30895 - 30899

  --0111100010110100    0111100010110101    0111100010110110    0111100010110111    0111100010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30900 - 30904

  --0111100010111001    0111100010111010    0111100010111011    0111100010111100    0111100010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30905 - 30909

  --0111100010111110    0111100010111111    0111100011000000    0111100011000001    0111100011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30910 - 30914

  --0111100011000011    0111100011000100    0111100011000101    0111100011000110    0111100011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30915 - 30919

  --0111100011001000    0111100011001001    0111100011001010    0111100011001011    0111100011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30920 - 30924

  --0111100011001101    0111100011001110    0111100011001111    0111100011010000    0111100011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30925 - 30929

  --0111100011010010    0111100011010011    0111100011010100    0111100011010101    0111100011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30930 - 30934

  --0111100011010111    0111100011011000    0111100011011001    0111100011011010    0111100011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30935 - 30939

  --0111100011011100    0111100011011101    0111100011011110    0111100011011111    0111100011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30940 - 30944

  --0111100011100001    0111100011100010    0111100011100011    0111100011100100    0111100011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30945 - 30949

  --0111100011100110    0111100011100111    0111100011101000    0111100011101001    0111100011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30950 - 30954

  --0111100011101011    0111100011101100    0111100011101101    0111100011101110    0111100011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30955 - 30959

  --0111100011110000    0111100011110001    0111100011110010    0111100011110011    0111100011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30960 - 30964

  --0111100011110101    0111100011110110    0111100011110111    0111100011111000    0111100011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30965 - 30969

  --0111100011111010    0111100011111011    0111100011111100    0111100011111101    0111100011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30970 - 30974

  --0111100011111111    0111100100000000    0111100100000001    0111100100000010    0111100100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30975 - 30979

  --0111100100000100    0111100100000101    0111100100000110    0111100100000111    0111100100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30980 - 30984

  --0111100100001001    0111100100001010    0111100100001011    0111100100001100    0111100100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30985 - 30989

  --0111100100001110    0111100100001111    0111100100010000    0111100100010001    0111100100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30990 - 30994

  --0111100100010011    0111100100010100    0111100100010101    0111100100010110    0111100100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 30995 - 30999

  --0111100100011000    0111100100011001    0111100100011010    0111100100011011    0111100100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31000 - 31004

  --0111100100011101    0111100100011110    0111100100011111    0111100100100000    0111100100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31005 - 31009

  --0111100100100010    0111100100100011    0111100100100100    0111100100100101    0111100100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31010 - 31014

  --0111100100100111    0111100100101000    0111100100101001    0111100100101010    0111100100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31015 - 31019

  --0111100100101100    0111100100101101    0111100100101110    0111100100101111    0111100100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31020 - 31024

  --0111100100110001    0111100100110010    0111100100110011    0111100100110100    0111100100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31025 - 31029

  --0111100100110110    0111100100110111    0111100100111000    0111100100111001    0111100100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31030 - 31034

  --0111100100111011    0111100100111100    0111100100111101    0111100100111110    0111100100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31035 - 31039

  --0111100101000000    0111100101000001    0111100101000010    0111100101000011    0111100101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31040 - 31044

  --0111100101000101    0111100101000110    0111100101000111    0111100101001000    0111100101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31045 - 31049

  --0111100101001010    0111100101001011    0111100101001100    0111100101001101    0111100101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31050 - 31054

  --0111100101001111    0111100101010000    0111100101010001    0111100101010010    0111100101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31055 - 31059

  --0111100101010100    0111100101010101    0111100101010110    0111100101010111    0111100101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31060 - 31064

  --0111100101011001    0111100101011010    0111100101011011    0111100101011100    0111100101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31065 - 31069

  --0111100101011110    0111100101011111    0111100101100000    0111100101100001    0111100101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31070 - 31074

  --0111100101100011    0111100101100100    0111100101100101    0111100101100110    0111100101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31075 - 31079

  --0111100101101000    0111100101101001    0111100101101010    0111100101101011    0111100101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31080 - 31084

  --0111100101101101    0111100101101110    0111100101101111    0111100101110000    0111100101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31085 - 31089

  --0111100101110010    0111100101110011    0111100101110100    0111100101110101    0111100101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31090 - 31094

  --0111100101110111    0111100101111000    0111100101111001    0111100101111010    0111100101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31095 - 31099

  --0111100101111100    0111100101111101    0111100101111110    0111100101111111    0111100110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31100 - 31104

  --0111100110000001    0111100110000010    0111100110000011    0111100110000100    0111100110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31105 - 31109

  --0111100110000110    0111100110000111    0111100110001000    0111100110001001    0111100110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31110 - 31114

  --0111100110001011    0111100110001100    0111100110001101    0111100110001110    0111100110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31115 - 31119

  --0111100110010000    0111100110010001    0111100110010010    0111100110010011    0111100110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31120 - 31124

  --0111100110010101    0111100110010110    0111100110010111    0111100110011000    0111100110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31125 - 31129

  --0111100110011010    0111100110011011    0111100110011100    0111100110011101    0111100110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31130 - 31134

  --0111100110011111    0111100110100000    0111100110100001    0111100110100010    0111100110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31135 - 31139

  --0111100110100100    0111100110100101    0111100110100110    0111100110100111    0111100110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31140 - 31144

  --0111100110101001    0111100110101010    0111100110101011    0111100110101100    0111100110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31145 - 31149

  --0111100110101110    0111100110101111    0111100110110000    0111100110110001    0111100110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31150 - 31154

  --0111100110110011    0111100110110100    0111100110110101    0111100110110110    0111100110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31155 - 31159

  --0111100110111000    0111100110111001    0111100110111010    0111100110111011    0111100110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31160 - 31164

  --0111100110111101    0111100110111110    0111100110111111    0111100111000000    0111100111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31165 - 31169

  --0111100111000010    0111100111000011    0111100111000100    0111100111000101    0111100111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31170 - 31174

  --0111100111000111    0111100111001000    0111100111001001    0111100111001010    0111100111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31175 - 31179

  --0111100111001100    0111100111001101    0111100111001110    0111100111001111    0111100111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31180 - 31184

  --0111100111010001    0111100111010010    0111100111010011    0111100111010100    0111100111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31185 - 31189

  --0111100111010110    0111100111010111    0111100111011000    0111100111011001    0111100111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31190 - 31194

  --0111100111011011    0111100111011100    0111100111011101    0111100111011110    0111100111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31195 - 31199

  --0111100111100000    0111100111100001    0111100111100010    0111100111100011    0111100111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31200 - 31204

  --0111100111100101    0111100111100110    0111100111100111    0111100111101000    0111100111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31205 - 31209

  --0111100111101010    0111100111101011    0111100111101100    0111100111101101    0111100111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31210 - 31214

  --0111100111101111    0111100111110000    0111100111110001    0111100111110010    0111100111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31215 - 31219

  --0111100111110100    0111100111110101    0111100111110110    0111100111110111    0111100111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31220 - 31224

  --0111100111111001    0111100111111010    0111100111111011    0111100111111100    0111100111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31225 - 31229

  --0111100111111110    0111100111111111    0111101000000000    0111101000000001    0111101000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31230 - 31234

  --0111101000000011    0111101000000100    0111101000000101    0111101000000110    0111101000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31235 - 31239

  --0111101000001000    0111101000001001    0111101000001010    0111101000001011    0111101000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31240 - 31244

  --0111101000001101    0111101000001110    0111101000001111    0111101000010000    0111101000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31245 - 31249

  --0111101000010010    0111101000010011    0111101000010100    0111101000010101    0111101000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31250 - 31254

  --0111101000010111    0111101000011000    0111101000011001    0111101000011010    0111101000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31255 - 31259

  --0111101000011100    0111101000011101    0111101000011110    0111101000011111    0111101000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31260 - 31264

  --0111101000100001    0111101000100010    0111101000100011    0111101000100100    0111101000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31265 - 31269

  --0111101000100110    0111101000100111    0111101000101000    0111101000101001    0111101000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31270 - 31274

  --0111101000101011    0111101000101100    0111101000101101    0111101000101110    0111101000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31275 - 31279

  --0111101000110000    0111101000110001    0111101000110010    0111101000110011    0111101000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31280 - 31284

  --0111101000110101    0111101000110110    0111101000110111    0111101000111000    0111101000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31285 - 31289

  --0111101000111010    0111101000111011    0111101000111100    0111101000111101    0111101000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31290 - 31294

  --0111101000111111    0111101001000000    0111101001000001    0111101001000010    0111101001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31295 - 31299

  --0111101001000100    0111101001000101    0111101001000110    0111101001000111    0111101001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31300 - 31304

  --0111101001001001    0111101001001010    0111101001001011    0111101001001100    0111101001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31305 - 31309

  --0111101001001110    0111101001001111    0111101001010000    0111101001010001    0111101001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31310 - 31314

  --0111101001010011    0111101001010100    0111101001010101    0111101001010110    0111101001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31315 - 31319

  --0111101001011000    0111101001011001    0111101001011010    0111101001011011    0111101001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31320 - 31324

  --0111101001011101    0111101001011110    0111101001011111    0111101001100000    0111101001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31325 - 31329

  --0111101001100010    0111101001100011    0111101001100100    0111101001100101    0111101001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31330 - 31334

  --0111101001100111    0111101001101000    0111101001101001    0111101001101010    0111101001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31335 - 31339

  --0111101001101100    0111101001101101    0111101001101110    0111101001101111    0111101001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31340 - 31344

  --0111101001110001    0111101001110010    0111101001110011    0111101001110100    0111101001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31345 - 31349

  --0111101001110110    0111101001110111    0111101001111000    0111101001111001    0111101001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31350 - 31354

  --0111101001111011    0111101001111100    0111101001111101    0111101001111110    0111101001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31355 - 31359

  --0111101010000000    0111101010000001    0111101010000010    0111101010000011    0111101010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31360 - 31364

  --0111101010000101    0111101010000110    0111101010000111    0111101010001000    0111101010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31365 - 31369

  --0111101010001010    0111101010001011    0111101010001100    0111101010001101    0111101010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31370 - 31374

  --0111101010001111    0111101010010000    0111101010010001    0111101010010010    0111101010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31375 - 31379

  --0111101010010100    0111101010010101    0111101010010110    0111101010010111    0111101010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31380 - 31384

  --0111101010011001    0111101010011010    0111101010011011    0111101010011100    0111101010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31385 - 31389

  --0111101010011110    0111101010011111    0111101010100000    0111101010100001    0111101010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31390 - 31394

  --0111101010100011    0111101010100100    0111101010100101    0111101010100110    0111101010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31395 - 31399

  --0111101010101000    0111101010101001    0111101010101010    0111101010101011    0111101010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31400 - 31404

  --0111101010101101    0111101010101110    0111101010101111    0111101010110000    0111101010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31405 - 31409

  --0111101010110010    0111101010110011    0111101010110100    0111101010110101    0111101010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31410 - 31414

  --0111101010110111    0111101010111000    0111101010111001    0111101010111010    0111101010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31415 - 31419

  --0111101010111100    0111101010111101    0111101010111110    0111101010111111    0111101011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31420 - 31424

  --0111101011000001    0111101011000010    0111101011000011    0111101011000100    0111101011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31425 - 31429

  --0111101011000110    0111101011000111    0111101011001000    0111101011001001    0111101011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31430 - 31434

  --0111101011001011    0111101011001100    0111101011001101    0111101011001110    0111101011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31435 - 31439

  --0111101011010000    0111101011010001    0111101011010010    0111101011010011    0111101011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31440 - 31444

  --0111101011010101    0111101011010110    0111101011010111    0111101011011000    0111101011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31445 - 31449

  --0111101011011010    0111101011011011    0111101011011100    0111101011011101    0111101011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31450 - 31454

  --0111101011011111    0111101011100000    0111101011100001    0111101011100010    0111101011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31455 - 31459

  --0111101011100100    0111101011100101    0111101011100110    0111101011100111    0111101011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31460 - 31464

  --0111101011101001    0111101011101010    0111101011101011    0111101011101100    0111101011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31465 - 31469

  --0111101011101110    0111101011101111    0111101011110000    0111101011110001    0111101011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31470 - 31474

  --0111101011110011    0111101011110100    0111101011110101    0111101011110110    0111101011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31475 - 31479

  --0111101011111000    0111101011111001    0111101011111010    0111101011111011    0111101011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31480 - 31484

  --0111101011111101    0111101011111110    0111101011111111    0111101100000000    0111101100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31485 - 31489

  --0111101100000010    0111101100000011    0111101100000100    0111101100000101    0111101100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31490 - 31494

  --0111101100000111    0111101100001000    0111101100001001    0111101100001010    0111101100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31495 - 31499

  --0111101100001100    0111101100001101    0111101100001110    0111101100001111    0111101100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31500 - 31504

  --0111101100010001    0111101100010010    0111101100010011    0111101100010100    0111101100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31505 - 31509

  --0111101100010110    0111101100010111    0111101100011000    0111101100011001    0111101100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31510 - 31514

  --0111101100011011    0111101100011100    0111101100011101    0111101100011110    0111101100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31515 - 31519

  --0111101100100000    0111101100100001    0111101100100010    0111101100100011    0111101100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31520 - 31524

  --0111101100100101    0111101100100110    0111101100100111    0111101100101000    0111101100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31525 - 31529

  --0111101100101010    0111101100101011    0111101100101100    0111101100101101    0111101100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31530 - 31534

  --0111101100101111    0111101100110000    0111101100110001    0111101100110010    0111101100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31535 - 31539

  --0111101100110100    0111101100110101    0111101100110110    0111101100110111    0111101100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31540 - 31544

  --0111101100111001    0111101100111010    0111101100111011    0111101100111100    0111101100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31545 - 31549

  --0111101100111110    0111101100111111    0111101101000000    0111101101000001    0111101101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31550 - 31554

  --0111101101000011    0111101101000100    0111101101000101    0111101101000110    0111101101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31555 - 31559

  --0111101101001000    0111101101001001    0111101101001010    0111101101001011    0111101101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31560 - 31564

  --0111101101001101    0111101101001110    0111101101001111    0111101101010000    0111101101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31565 - 31569

  --0111101101010010    0111101101010011    0111101101010100    0111101101010101    0111101101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31570 - 31574

  --0111101101010111    0111101101011000    0111101101011001    0111101101011010    0111101101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31575 - 31579

  --0111101101011100    0111101101011101    0111101101011110    0111101101011111    0111101101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31580 - 31584

  --0111101101100001    0111101101100010    0111101101100011    0111101101100100    0111101101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31585 - 31589

  --0111101101100110    0111101101100111    0111101101101000    0111101101101001    0111101101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31590 - 31594

  --0111101101101011    0111101101101100    0111101101101101    0111101101101110    0111101101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31595 - 31599

  --0111101101110000    0111101101110001    0111101101110010    0111101101110011    0111101101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31600 - 31604

  --0111101101110101    0111101101110110    0111101101110111    0111101101111000    0111101101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31605 - 31609

  --0111101101111010    0111101101111011    0111101101111100    0111101101111101    0111101101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31610 - 31614

  --0111101101111111    0111101110000000    0111101110000001    0111101110000010    0111101110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31615 - 31619

  --0111101110000100    0111101110000101    0111101110000110    0111101110000111    0111101110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31620 - 31624

  --0111101110001001    0111101110001010    0111101110001011    0111101110001100    0111101110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31625 - 31629

  --0111101110001110    0111101110001111    0111101110010000    0111101110010001    0111101110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31630 - 31634

  --0111101110010011    0111101110010100    0111101110010101    0111101110010110    0111101110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31635 - 31639

  --0111101110011000    0111101110011001    0111101110011010    0111101110011011    0111101110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31640 - 31644

  --0111101110011101    0111101110011110    0111101110011111    0111101110100000    0111101110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31645 - 31649

  --0111101110100010    0111101110100011    0111101110100100    0111101110100101    0111101110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31650 - 31654

  --0111101110100111    0111101110101000    0111101110101001    0111101110101010    0111101110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31655 - 31659

  --0111101110101100    0111101110101101    0111101110101110    0111101110101111    0111101110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31660 - 31664

  --0111101110110001    0111101110110010    0111101110110011    0111101110110100    0111101110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31665 - 31669

  --0111101110110110    0111101110110111    0111101110111000    0111101110111001    0111101110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31670 - 31674

  --0111101110111011    0111101110111100    0111101110111101    0111101110111110    0111101110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31675 - 31679

  --0111101111000000    0111101111000001    0111101111000010    0111101111000011    0111101111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31680 - 31684

  --0111101111000101    0111101111000110    0111101111000111    0111101111001000    0111101111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31685 - 31689

  --0111101111001010    0111101111001011    0111101111001100    0111101111001101    0111101111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31690 - 31694

  --0111101111001111    0111101111010000    0111101111010001    0111101111010010    0111101111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31695 - 31699

  --0111101111010100    0111101111010101    0111101111010110    0111101111010111    0111101111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31700 - 31704

  --0111101111011001    0111101111011010    0111101111011011    0111101111011100    0111101111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31705 - 31709

  --0111101111011110    0111101111011111    0111101111100000    0111101111100001    0111101111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31710 - 31714

  --0111101111100011    0111101111100100    0111101111100101    0111101111100110    0111101111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31715 - 31719

  --0111101111101000    0111101111101001    0111101111101010    0111101111101011    0111101111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31720 - 31724

  --0111101111101101    0111101111101110    0111101111101111    0111101111110000    0111101111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31725 - 31729

  --0111101111110010    0111101111110011    0111101111110100    0111101111110101    0111101111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31730 - 31734

  --0111101111110111    0111101111111000    0111101111111001    0111101111111010    0111101111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31735 - 31739

  --0111101111111100    0111101111111101    0111101111111110    0111101111111111    0111110000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31740 - 31744

  --0111110000000001    0111110000000010    0111110000000011    0111110000000100    0111110000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31745 - 31749

  --0111110000000110    0111110000000111    0111110000001000    0111110000001001    0111110000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31750 - 31754

  --0111110000001011    0111110000001100    0111110000001101    0111110000001110    0111110000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31755 - 31759

  --0111110000010000    0111110000010001    0111110000010010    0111110000010011    0111110000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31760 - 31764

  --0111110000010101    0111110000010110    0111110000010111    0111110000011000    0111110000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31765 - 31769

  --0111110000011010    0111110000011011    0111110000011100    0111110000011101    0111110000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31770 - 31774

  --0111110000011111    0111110000100000    0111110000100001    0111110000100010    0111110000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31775 - 31779

  --0111110000100100    0111110000100101    0111110000100110    0111110000100111    0111110000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31780 - 31784

  --0111110000101001    0111110000101010    0111110000101011    0111110000101100    0111110000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31785 - 31789

  --0111110000101110    0111110000101111    0111110000110000    0111110000110001    0111110000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31790 - 31794

  --0111110000110011    0111110000110100    0111110000110101    0111110000110110    0111110000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31795 - 31799

  --0111110000111000    0111110000111001    0111110000111010    0111110000111011    0111110000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31800 - 31804

  --0111110000111101    0111110000111110    0111110000111111    0111110001000000    0111110001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31805 - 31809

  --0111110001000010    0111110001000011    0111110001000100    0111110001000101    0111110001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31810 - 31814

  --0111110001000111    0111110001001000    0111110001001001    0111110001001010    0111110001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31815 - 31819

  --0111110001001100    0111110001001101    0111110001001110    0111110001001111    0111110001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31820 - 31824

  --0111110001010001    0111110001010010    0111110001010011    0111110001010100    0111110001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31825 - 31829

  --0111110001010110    0111110001010111    0111110001011000    0111110001011001    0111110001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31830 - 31834

  --0111110001011011    0111110001011100    0111110001011101    0111110001011110    0111110001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31835 - 31839

  --0111110001100000    0111110001100001    0111110001100010    0111110001100011    0111110001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31840 - 31844

  --0111110001100101    0111110001100110    0111110001100111    0111110001101000    0111110001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31845 - 31849

  --0111110001101010    0111110001101011    0111110001101100    0111110001101101    0111110001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31850 - 31854

  --0111110001101111    0111110001110000    0111110001110001    0111110001110010    0111110001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31855 - 31859

  --0111110001110100    0111110001110101    0111110001110110    0111110001110111    0111110001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31860 - 31864

  --0111110001111001    0111110001111010    0111110001111011    0111110001111100    0111110001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31865 - 31869

  --0111110001111110    0111110001111111    0111110010000000    0111110010000001    0111110010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31870 - 31874

  --0111110010000011    0111110010000100    0111110010000101    0111110010000110    0111110010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31875 - 31879

  --0111110010001000    0111110010001001    0111110010001010    0111110010001011    0111110010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31880 - 31884

  --0111110010001101    0111110010001110    0111110010001111    0111110010010000    0111110010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31885 - 31889

  --0111110010010010    0111110010010011    0111110010010100    0111110010010101    0111110010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31890 - 31894

  --0111110010010111    0111110010011000    0111110010011001    0111110010011010    0111110010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31895 - 31899

  --0111110010011100    0111110010011101    0111110010011110    0111110010011111    0111110010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31900 - 31904

  --0111110010100001    0111110010100010    0111110010100011    0111110010100100    0111110010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31905 - 31909

  --0111110010100110    0111110010100111    0111110010101000    0111110010101001    0111110010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31910 - 31914

  --0111110010101011    0111110010101100    0111110010101101    0111110010101110    0111110010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31915 - 31919

  --0111110010110000    0111110010110001    0111110010110010    0111110010110011    0111110010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31920 - 31924

  --0111110010110101    0111110010110110    0111110010110111    0111110010111000    0111110010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31925 - 31929

  --0111110010111010    0111110010111011    0111110010111100    0111110010111101    0111110010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31930 - 31934

  --0111110010111111    0111110011000000    0111110011000001    0111110011000010    0111110011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31935 - 31939

  --0111110011000100    0111110011000101    0111110011000110    0111110011000111    0111110011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31940 - 31944

  --0111110011001001    0111110011001010    0111110011001011    0111110011001100    0111110011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31945 - 31949

  --0111110011001110    0111110011001111    0111110011010000    0111110011010001    0111110011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31950 - 31954

  --0111110011010011    0111110011010100    0111110011010101    0111110011010110    0111110011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31955 - 31959

  --0111110011011000    0111110011011001    0111110011011010    0111110011011011    0111110011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31960 - 31964

  --0111110011011101    0111110011011110    0111110011011111    0111110011100000    0111110011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31965 - 31969

  --0111110011100010    0111110011100011    0111110011100100    0111110011100101    0111110011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31970 - 31974

  --0111110011100111    0111110011101000    0111110011101001    0111110011101010    0111110011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31975 - 31979

  --0111110011101100    0111110011101101    0111110011101110    0111110011101111    0111110011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31980 - 31984

  --0111110011110001    0111110011110010    0111110011110011    0111110011110100    0111110011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31985 - 31989

  --0111110011110110    0111110011110111    0111110011111000    0111110011111001    0111110011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31990 - 31994

  --0111110011111011    0111110011111100    0111110011111101    0111110011111110    0111110011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 31995 - 31999

  --0111110100000000    0111110100000001    0111110100000010    0111110100000011    0111110100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32000 - 32004

  --0111110100000101    0111110100000110    0111110100000111    0111110100001000    0111110100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32005 - 32009

  --0111110100001010    0111110100001011    0111110100001100    0111110100001101    0111110100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32010 - 32014

  --0111110100001111    0111110100010000    0111110100010001    0111110100010010    0111110100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32015 - 32019

  --0111110100010100    0111110100010101    0111110100010110    0111110100010111    0111110100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32020 - 32024

  --0111110100011001    0111110100011010    0111110100011011    0111110100011100    0111110100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32025 - 32029

  --0111110100011110    0111110100011111    0111110100100000    0111110100100001    0111110100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32030 - 32034

  --0111110100100011    0111110100100100    0111110100100101    0111110100100110    0111110100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32035 - 32039

  --0111110100101000    0111110100101001    0111110100101010    0111110100101011    0111110100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32040 - 32044

  --0111110100101101    0111110100101110    0111110100101111    0111110100110000    0111110100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32045 - 32049

  --0111110100110010    0111110100110011    0111110100110100    0111110100110101    0111110100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32050 - 32054

  --0111110100110111    0111110100111000    0111110100111001    0111110100111010    0111110100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32055 - 32059

  --0111110100111100    0111110100111101    0111110100111110    0111110100111111    0111110101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32060 - 32064

  --0111110101000001    0111110101000010    0111110101000011    0111110101000100    0111110101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32065 - 32069

  --0111110101000110    0111110101000111    0111110101001000    0111110101001001    0111110101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32070 - 32074

  --0111110101001011    0111110101001100    0111110101001101    0111110101001110    0111110101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32075 - 32079

  --0111110101010000    0111110101010001    0111110101010010    0111110101010011    0111110101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32080 - 32084

  --0111110101010101    0111110101010110    0111110101010111    0111110101011000    0111110101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32085 - 32089

  --0111110101011010    0111110101011011    0111110101011100    0111110101011101    0111110101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32090 - 32094

  --0111110101011111    0111110101100000    0111110101100001    0111110101100010    0111110101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32095 - 32099

  --0111110101100100    0111110101100101    0111110101100110    0111110101100111    0111110101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32100 - 32104

  --0111110101101001    0111110101101010    0111110101101011    0111110101101100    0111110101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32105 - 32109

  --0111110101101110    0111110101101111    0111110101110000    0111110101110001    0111110101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32110 - 32114

  --0111110101110011    0111110101110100    0111110101110101    0111110101110110    0111110101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32115 - 32119

  --0111110101111000    0111110101111001    0111110101111010    0111110101111011    0111110101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32120 - 32124

  --0111110101111101    0111110101111110    0111110101111111    0111110110000000    0111110110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32125 - 32129

  --0111110110000010    0111110110000011    0111110110000100    0111110110000101    0111110110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32130 - 32134

  --0111110110000111    0111110110001000    0111110110001001    0111110110001010    0111110110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32135 - 32139

  --0111110110001100    0111110110001101    0111110110001110    0111110110001111    0111110110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32140 - 32144

  --0111110110010001    0111110110010010    0111110110010011    0111110110010100    0111110110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32145 - 32149

  --0111110110010110    0111110110010111    0111110110011000    0111110110011001    0111110110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32150 - 32154

  --0111110110011011    0111110110011100    0111110110011101    0111110110011110    0111110110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32155 - 32159

  --0111110110100000    0111110110100001    0111110110100010    0111110110100011    0111110110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32160 - 32164

  --0111110110100101    0111110110100110    0111110110100111    0111110110101000    0111110110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32165 - 32169

  --0111110110101010    0111110110101011    0111110110101100    0111110110101101    0111110110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32170 - 32174

  --0111110110101111    0111110110110000    0111110110110001    0111110110110010    0111110110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32175 - 32179

  --0111110110110100    0111110110110101    0111110110110110    0111110110110111    0111110110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32180 - 32184

  --0111110110111001    0111110110111010    0111110110111011    0111110110111100    0111110110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32185 - 32189

  --0111110110111110    0111110110111111    0111110111000000    0111110111000001    0111110111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32190 - 32194

  --0111110111000011    0111110111000100    0111110111000101    0111110111000110    0111110111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32195 - 32199

  --0111110111001000    0111110111001001    0111110111001010    0111110111001011    0111110111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32200 - 32204

  --0111110111001101    0111110111001110    0111110111001111    0111110111010000    0111110111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32205 - 32209

  --0111110111010010    0111110111010011    0111110111010100    0111110111010101    0111110111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32210 - 32214

  --0111110111010111    0111110111011000    0111110111011001    0111110111011010    0111110111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32215 - 32219

  --0111110111011100    0111110111011101    0111110111011110    0111110111011111    0111110111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32220 - 32224

  --0111110111100001    0111110111100010    0111110111100011    0111110111100100    0111110111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32225 - 32229

  --0111110111100110    0111110111100111    0111110111101000    0111110111101001    0111110111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32230 - 32234

  --0111110111101011    0111110111101100    0111110111101101    0111110111101110    0111110111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32235 - 32239

  --0111110111110000    0111110111110001    0111110111110010    0111110111110011    0111110111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32240 - 32244

  --0111110111110101    0111110111110110    0111110111110111    0111110111111000    0111110111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32245 - 32249

  --0111110111111010    0111110111111011    0111110111111100    0111110111111101    0111110111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32250 - 32254

  --0111110111111111    0111111000000000    0111111000000001    0111111000000010    0111111000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32255 - 32259

  --0111111000000100    0111111000000101    0111111000000110    0111111000000111    0111111000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32260 - 32264

  --0111111000001001    0111111000001010    0111111000001011    0111111000001100    0111111000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32265 - 32269

  --0111111000001110    0111111000001111    0111111000010000    0111111000010001    0111111000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32270 - 32274

  --0111111000010011    0111111000010100    0111111000010101    0111111000010110    0111111000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32275 - 32279

  --0111111000011000    0111111000011001    0111111000011010    0111111000011011    0111111000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32280 - 32284

  --0111111000011101    0111111000011110    0111111000011111    0111111000100000    0111111000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32285 - 32289

  --0111111000100010    0111111000100011    0111111000100100    0111111000100101    0111111000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32290 - 32294

  --0111111000100111    0111111000101000    0111111000101001    0111111000101010    0111111000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32295 - 32299

  --0111111000101100    0111111000101101    0111111000101110    0111111000101111    0111111000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32300 - 32304

  --0111111000110001    0111111000110010    0111111000110011    0111111000110100    0111111000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32305 - 32309

  --0111111000110110    0111111000110111    0111111000111000    0111111000111001    0111111000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32310 - 32314

  --0111111000111011    0111111000111100    0111111000111101    0111111000111110    0111111000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32315 - 32319

  --0111111001000000    0111111001000001    0111111001000010    0111111001000011    0111111001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32320 - 32324

  --0111111001000101    0111111001000110    0111111001000111    0111111001001000    0111111001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32325 - 32329

  --0111111001001010    0111111001001011    0111111001001100    0111111001001101    0111111001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32330 - 32334

  --0111111001001111    0111111001010000    0111111001010001    0111111001010010    0111111001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32335 - 32339

  --0111111001010100    0111111001010101    0111111001010110    0111111001010111    0111111001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32340 - 32344

  --0111111001011001    0111111001011010    0111111001011011    0111111001011100    0111111001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32345 - 32349

  --0111111001011110    0111111001011111    0111111001100000    0111111001100001    0111111001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32350 - 32354

  --0111111001100011    0111111001100100    0111111001100101    0111111001100110    0111111001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32355 - 32359

  --0111111001101000    0111111001101001    0111111001101010    0111111001101011    0111111001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32360 - 32364

  --0111111001101101    0111111001101110    0111111001101111    0111111001110000    0111111001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32365 - 32369

  --0111111001110010    0111111001110011    0111111001110100    0111111001110101    0111111001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32370 - 32374

  --0111111001110111    0111111001111000    0111111001111001    0111111001111010    0111111001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32375 - 32379

  --0111111001111100    0111111001111101    0111111001111110    0111111001111111    0111111010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32380 - 32384

  --0111111010000001    0111111010000010    0111111010000011    0111111010000100    0111111010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32385 - 32389

  --0111111010000110    0111111010000111    0111111010001000    0111111010001001    0111111010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32390 - 32394

  --0111111010001011    0111111010001100    0111111010001101    0111111010001110    0111111010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32395 - 32399

  --0111111010010000    0111111010010001    0111111010010010    0111111010010011    0111111010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32400 - 32404

  --0111111010010101    0111111010010110    0111111010010111    0111111010011000    0111111010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32405 - 32409

  --0111111010011010    0111111010011011    0111111010011100    0111111010011101    0111111010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32410 - 32414

  --0111111010011111    0111111010100000    0111111010100001    0111111010100010    0111111010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32415 - 32419

  --0111111010100100    0111111010100101    0111111010100110    0111111010100111    0111111010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32420 - 32424

  --0111111010101001    0111111010101010    0111111010101011    0111111010101100    0111111010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32425 - 32429

  --0111111010101110    0111111010101111    0111111010110000    0111111010110001    0111111010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32430 - 32434

  --0111111010110011    0111111010110100    0111111010110101    0111111010110110    0111111010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32435 - 32439

  --0111111010111000    0111111010111001    0111111010111010    0111111010111011    0111111010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32440 - 32444

  --0111111010111101    0111111010111110    0111111010111111    0111111011000000    0111111011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32445 - 32449

  --0111111011000010    0111111011000011    0111111011000100    0111111011000101    0111111011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32450 - 32454

  --0111111011000111    0111111011001000    0111111011001001    0111111011001010    0111111011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32455 - 32459

  --0111111011001100    0111111011001101    0111111011001110    0111111011001111    0111111011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32460 - 32464

  --0111111011010001    0111111011010010    0111111011010011    0111111011010100    0111111011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32465 - 32469

  --0111111011010110    0111111011010111    0111111011011000    0111111011011001    0111111011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32470 - 32474

  --0111111011011011    0111111011011100    0111111011011101    0111111011011110    0111111011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32475 - 32479

  --0111111011100000    0111111011100001    0111111011100010    0111111011100011    0111111011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32480 - 32484

  --0111111011100101    0111111011100110    0111111011100111    0111111011101000    0111111011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32485 - 32489

  --0111111011101010    0111111011101011    0111111011101100    0111111011101101    0111111011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32490 - 32494

  --0111111011101111    0111111011110000    0111111011110001    0111111011110010    0111111011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32495 - 32499

  --0111111011110100    0111111011110101    0111111011110110    0111111011110111    0111111011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32500 - 32504

  --0111111011111001    0111111011111010    0111111011111011    0111111011111100    0111111011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32505 - 32509

  --0111111011111110    0111111011111111    0111111100000000    0111111100000001    0111111100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32510 - 32514

  --0111111100000011    0111111100000100    0111111100000101    0111111100000110    0111111100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32515 - 32519

  --0111111100001000    0111111100001001    0111111100001010    0111111100001011    0111111100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32520 - 32524

  --0111111100001101    0111111100001110    0111111100001111    0111111100010000    0111111100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32525 - 32529

  --0111111100010010    0111111100010011    0111111100010100    0111111100010101    0111111100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32530 - 32534

  --0111111100010111    0111111100011000    0111111100011001    0111111100011010    0111111100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32535 - 32539

  --0111111100011100    0111111100011101    0111111100011110    0111111100011111    0111111100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32540 - 32544

  --0111111100100001    0111111100100010    0111111100100011    0111111100100100    0111111100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32545 - 32549

  --0111111100100110    0111111100100111    0111111100101000    0111111100101001    0111111100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32550 - 32554

  --0111111100101011    0111111100101100    0111111100101101    0111111100101110    0111111100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32555 - 32559

  --0111111100110000    0111111100110001    0111111100110010    0111111100110011    0111111100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32560 - 32564

  --0111111100110101    0111111100110110    0111111100110111    0111111100111000    0111111100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32565 - 32569

  --0111111100111010    0111111100111011    0111111100111100    0111111100111101    0111111100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32570 - 32574

  --0111111100111111    0111111101000000    0111111101000001    0111111101000010    0111111101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32575 - 32579

  --0111111101000100    0111111101000101    0111111101000110    0111111101000111    0111111101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32580 - 32584

  --0111111101001001    0111111101001010    0111111101001011    0111111101001100    0111111101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32585 - 32589

  --0111111101001110    0111111101001111    0111111101010000    0111111101010001    0111111101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32590 - 32594

  --0111111101010011    0111111101010100    0111111101010101    0111111101010110    0111111101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32595 - 32599

  --0111111101011000    0111111101011001    0111111101011010    0111111101011011    0111111101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32600 - 32604

  --0111111101011101    0111111101011110    0111111101011111    0111111101100000    0111111101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32605 - 32609

  --0111111101100010    0111111101100011    0111111101100100    0111111101100101    0111111101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32610 - 32614

  --0111111101100111    0111111101101000    0111111101101001    0111111101101010    0111111101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32615 - 32619

  --0111111101101100    0111111101101101    0111111101101110    0111111101101111    0111111101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32620 - 32624

  --0111111101110001    0111111101110010    0111111101110011    0111111101110100    0111111101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32625 - 32629

  --0111111101110110    0111111101110111    0111111101111000    0111111101111001    0111111101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32630 - 32634

  --0111111101111011    0111111101111100    0111111101111101    0111111101111110    0111111101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32635 - 32639

  --0111111110000000    0111111110000001    0111111110000010    0111111110000011    0111111110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32640 - 32644

  --0111111110000101    0111111110000110    0111111110000111    0111111110001000    0111111110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32645 - 32649

  --0111111110001010    0111111110001011    0111111110001100    0111111110001101    0111111110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32650 - 32654

  --0111111110001111    0111111110010000    0111111110010001    0111111110010010    0111111110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32655 - 32659

  --0111111110010100    0111111110010101    0111111110010110    0111111110010111    0111111110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32660 - 32664

  --0111111110011001    0111111110011010    0111111110011011    0111111110011100    0111111110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32665 - 32669

  --0111111110011110    0111111110011111    0111111110100000    0111111110100001    0111111110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32670 - 32674

  --0111111110100011    0111111110100100    0111111110100101    0111111110100110    0111111110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32675 - 32679

  --0111111110101000    0111111110101001    0111111110101010    0111111110101011    0111111110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32680 - 32684

  --0111111110101101    0111111110101110    0111111110101111    0111111110110000    0111111110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32685 - 32689

  --0111111110110010    0111111110110011    0111111110110100    0111111110110101    0111111110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32690 - 32694

  --0111111110110111    0111111110111000    0111111110111001    0111111110111010    0111111110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32695 - 32699

  --0111111110111100    0111111110111101    0111111110111110    0111111110111111    0111111111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32700 - 32704

  --0111111111000001    0111111111000010    0111111111000011    0111111111000100    0111111111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32705 - 32709

  --0111111111000110    0111111111000111    0111111111001000    0111111111001001    0111111111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32710 - 32714

  --0111111111001011    0111111111001100    0111111111001101    0111111111001110    0111111111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32715 - 32719

  --0111111111010000    0111111111010001    0111111111010010    0111111111010011    0111111111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32720 - 32724

  --0111111111010101    0111111111010110    0111111111010111    0111111111011000    0111111111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32725 - 32729

  --0111111111011010    0111111111011011    0111111111011100    0111111111011101    0111111111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32730 - 32734

  --0111111111011111    0111111111100000    0111111111100001    0111111111100010    0111111111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32735 - 32739

  --0111111111100100    0111111111100101    0111111111100110    0111111111100111    0111111111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32740 - 32744

  --0111111111101001    0111111111101010    0111111111101011    0111111111101100    0111111111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32745 - 32749

  --0111111111101110    0111111111101111    0111111111110000    0111111111110001    0111111111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32750 - 32754

  --0111111111110011    0111111111110100    0111111111110101    0111111111110110    0111111111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32755 - 32759

  --0111111111111000    0111111111111001    0111111111111010    0111111111111011    0111111111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32760 - 32764

  --0111111111111101    0111111111111110    0111111111111111    1000000000000000    1000000000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32765 - 32769

  --1000000000000010    1000000000000011    1000000000000100    1000000000000101    1000000000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32770 - 32774

  --1000000000000111    1000000000001000    1000000000001001    1000000000001010    1000000000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32775 - 32779

  --1000000000001100    1000000000001101    1000000000001110    1000000000001111    1000000000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32780 - 32784

  --1000000000010001    1000000000010010    1000000000010011    1000000000010100    1000000000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32785 - 32789

  --1000000000010110    1000000000010111    1000000000011000    1000000000011001    1000000000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32790 - 32794

  --1000000000011011    1000000000011100    1000000000011101    1000000000011110    1000000000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32795 - 32799

  --1000000000100000    1000000000100001    1000000000100010    1000000000100011    1000000000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32800 - 32804

  --1000000000100101    1000000000100110    1000000000100111    1000000000101000    1000000000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32805 - 32809

  --1000000000101010    1000000000101011    1000000000101100    1000000000101101    1000000000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32810 - 32814

  --1000000000101111    1000000000110000    1000000000110001    1000000000110010    1000000000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32815 - 32819

  --1000000000110100    1000000000110101    1000000000110110    1000000000110111    1000000000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32820 - 32824

  --1000000000111001    1000000000111010    1000000000111011    1000000000111100    1000000000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32825 - 32829

  --1000000000111110    1000000000111111    1000000001000000    1000000001000001    1000000001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32830 - 32834

  --1000000001000011    1000000001000100    1000000001000101    1000000001000110    1000000001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32835 - 32839

  --1000000001001000    1000000001001001    1000000001001010    1000000001001011    1000000001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32840 - 32844

  --1000000001001101    1000000001001110    1000000001001111    1000000001010000    1000000001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32845 - 32849

  --1000000001010010    1000000001010011    1000000001010100    1000000001010101    1000000001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32850 - 32854

  --1000000001010111    1000000001011000    1000000001011001    1000000001011010    1000000001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32855 - 32859

  --1000000001011100    1000000001011101    1000000001011110    1000000001011111    1000000001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32860 - 32864

  --1000000001100001    1000000001100010    1000000001100011    1000000001100100    1000000001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32865 - 32869

  --1000000001100110    1000000001100111    1000000001101000    1000000001101001    1000000001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32870 - 32874

  --1000000001101011    1000000001101100    1000000001101101    1000000001101110    1000000001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32875 - 32879

  --1000000001110000    1000000001110001    1000000001110010    1000000001110011    1000000001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32880 - 32884

  --1000000001110101    1000000001110110    1000000001110111    1000000001111000    1000000001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32885 - 32889

  --1000000001111010    1000000001111011    1000000001111100    1000000001111101    1000000001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32890 - 32894

  --1000000001111111    1000000010000000    1000000010000001    1000000010000010    1000000010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32895 - 32899

  --1000000010000100    1000000010000101    1000000010000110    1000000010000111    1000000010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32900 - 32904

  --1000000010001001    1000000010001010    1000000010001011    1000000010001100    1000000010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32905 - 32909

  --1000000010001110    1000000010001111    1000000010010000    1000000010010001    1000000010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32910 - 32914

  --1000000010010011    1000000010010100    1000000010010101    1000000010010110    1000000010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32915 - 32919

  --1000000010011000    1000000010011001    1000000010011010    1000000010011011    1000000010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32920 - 32924

  --1000000010011101    1000000010011110    1000000010011111    1000000010100000    1000000010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32925 - 32929

  --1000000010100010    1000000010100011    1000000010100100    1000000010100101    1000000010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32930 - 32934

  --1000000010100111    1000000010101000    1000000010101001    1000000010101010    1000000010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32935 - 32939

  --1000000010101100    1000000010101101    1000000010101110    1000000010101111    1000000010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32940 - 32944

  --1000000010110001    1000000010110010    1000000010110011    1000000010110100    1000000010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32945 - 32949

  --1000000010110110    1000000010110111    1000000010111000    1000000010111001    1000000010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32950 - 32954

  --1000000010111011    1000000010111100    1000000010111101    1000000010111110    1000000010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32955 - 32959

  --1000000011000000    1000000011000001    1000000011000010    1000000011000011    1000000011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32960 - 32964

  --1000000011000101    1000000011000110    1000000011000111    1000000011001000    1000000011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32965 - 32969

  --1000000011001010    1000000011001011    1000000011001100    1000000011001101    1000000011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32970 - 32974

  --1000000011001111    1000000011010000    1000000011010001    1000000011010010    1000000011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32975 - 32979

  --1000000011010100    1000000011010101    1000000011010110    1000000011010111    1000000011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32980 - 32984

  --1000000011011001    1000000011011010    1000000011011011    1000000011011100    1000000011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32985 - 32989

  --1000000011011110    1000000011011111    1000000011100000    1000000011100001    1000000011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32990 - 32994

  --1000000011100011    1000000011100100    1000000011100101    1000000011100110    1000000011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 32995 - 32999

  --1000000011101000    1000000011101001    1000000011101010    1000000011101011    1000000011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33000 - 33004

  --1000000011101101    1000000011101110    1000000011101111    1000000011110000    1000000011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33005 - 33009

  --1000000011110010    1000000011110011    1000000011110100    1000000011110101    1000000011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33010 - 33014

  --1000000011110111    1000000011111000    1000000011111001    1000000011111010    1000000011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33015 - 33019

  --1000000011111100    1000000011111101    1000000011111110    1000000011111111    1000000100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33020 - 33024

  --1000000100000001    1000000100000010    1000000100000011    1000000100000100    1000000100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33025 - 33029

  --1000000100000110    1000000100000111    1000000100001000    1000000100001001    1000000100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33030 - 33034

  --1000000100001011    1000000100001100    1000000100001101    1000000100001110    1000000100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33035 - 33039

  --1000000100010000    1000000100010001    1000000100010010    1000000100010011    1000000100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33040 - 33044

  --1000000100010101    1000000100010110    1000000100010111    1000000100011000    1000000100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33045 - 33049

  --1000000100011010    1000000100011011    1000000100011100    1000000100011101    1000000100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33050 - 33054

  --1000000100011111    1000000100100000    1000000100100001    1000000100100010    1000000100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33055 - 33059

  --1000000100100100    1000000100100101    1000000100100110    1000000100100111    1000000100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33060 - 33064

  --1000000100101001    1000000100101010    1000000100101011    1000000100101100    1000000100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33065 - 33069

  --1000000100101110    1000000100101111    1000000100110000    1000000100110001    1000000100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33070 - 33074

  --1000000100110011    1000000100110100    1000000100110101    1000000100110110    1000000100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33075 - 33079

  --1000000100111000    1000000100111001    1000000100111010    1000000100111011    1000000100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33080 - 33084

  --1000000100111101    1000000100111110    1000000100111111    1000000101000000    1000000101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33085 - 33089

  --1000000101000010    1000000101000011    1000000101000100    1000000101000101    1000000101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33090 - 33094

  --1000000101000111    1000000101001000    1000000101001001    1000000101001010    1000000101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33095 - 33099

  --1000000101001100    1000000101001101    1000000101001110    1000000101001111    1000000101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33100 - 33104

  --1000000101010001    1000000101010010    1000000101010011    1000000101010100    1000000101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33105 - 33109

  --1000000101010110    1000000101010111    1000000101011000    1000000101011001    1000000101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33110 - 33114

  --1000000101011011    1000000101011100    1000000101011101    1000000101011110    1000000101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33115 - 33119

  --1000000101100000    1000000101100001    1000000101100010    1000000101100011    1000000101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33120 - 33124

  --1000000101100101    1000000101100110    1000000101100111    1000000101101000    1000000101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33125 - 33129

  --1000000101101010    1000000101101011    1000000101101100    1000000101101101    1000000101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33130 - 33134

  --1000000101101111    1000000101110000    1000000101110001    1000000101110010    1000000101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33135 - 33139

  --1000000101110100    1000000101110101    1000000101110110    1000000101110111    1000000101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33140 - 33144

  --1000000101111001    1000000101111010    1000000101111011    1000000101111100    1000000101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33145 - 33149

  --1000000101111110    1000000101111111    1000000110000000    1000000110000001    1000000110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33150 - 33154

  --1000000110000011    1000000110000100    1000000110000101    1000000110000110    1000000110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33155 - 33159

  --1000000110001000    1000000110001001    1000000110001010    1000000110001011    1000000110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33160 - 33164

  --1000000110001101    1000000110001110    1000000110001111    1000000110010000    1000000110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33165 - 33169

  --1000000110010010    1000000110010011    1000000110010100    1000000110010101    1000000110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33170 - 33174

  --1000000110010111    1000000110011000    1000000110011001    1000000110011010    1000000110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33175 - 33179

  --1000000110011100    1000000110011101    1000000110011110    1000000110011111    1000000110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33180 - 33184

  --1000000110100001    1000000110100010    1000000110100011    1000000110100100    1000000110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33185 - 33189

  --1000000110100110    1000000110100111    1000000110101000    1000000110101001    1000000110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33190 - 33194

  --1000000110101011    1000000110101100    1000000110101101    1000000110101110    1000000110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33195 - 33199

  --1000000110110000    1000000110110001    1000000110110010    1000000110110011    1000000110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33200 - 33204

  --1000000110110101    1000000110110110    1000000110110111    1000000110111000    1000000110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33205 - 33209

  --1000000110111010    1000000110111011    1000000110111100    1000000110111101    1000000110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33210 - 33214

  --1000000110111111    1000000111000000    1000000111000001    1000000111000010    1000000111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33215 - 33219

  --1000000111000100    1000000111000101    1000000111000110    1000000111000111    1000000111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33220 - 33224

  --1000000111001001    1000000111001010    1000000111001011    1000000111001100    1000000111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33225 - 33229

  --1000000111001110    1000000111001111    1000000111010000    1000000111010001    1000000111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33230 - 33234

  --1000000111010011    1000000111010100    1000000111010101    1000000111010110    1000000111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33235 - 33239

  --1000000111011000    1000000111011001    1000000111011010    1000000111011011    1000000111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33240 - 33244

  --1000000111011101    1000000111011110    1000000111011111    1000000111100000    1000000111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33245 - 33249

  --1000000111100010    1000000111100011    1000000111100100    1000000111100101    1000000111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33250 - 33254

  --1000000111100111    1000000111101000    1000000111101001    1000000111101010    1000000111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33255 - 33259

  --1000000111101100    1000000111101101    1000000111101110    1000000111101111    1000000111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33260 - 33264

  --1000000111110001    1000000111110010    1000000111110011    1000000111110100    1000000111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33265 - 33269

  --1000000111110110    1000000111110111    1000000111111000    1000000111111001    1000000111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33270 - 33274

  --1000000111111011    1000000111111100    1000000111111101    1000000111111110    1000000111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33275 - 33279

  --1000001000000000    1000001000000001    1000001000000010    1000001000000011    1000001000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33280 - 33284

  --1000001000000101    1000001000000110    1000001000000111    1000001000001000    1000001000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33285 - 33289

  --1000001000001010    1000001000001011    1000001000001100    1000001000001101    1000001000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33290 - 33294

  --1000001000001111    1000001000010000    1000001000010001    1000001000010010    1000001000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33295 - 33299

  --1000001000010100    1000001000010101    1000001000010110    1000001000010111    1000001000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33300 - 33304

  --1000001000011001    1000001000011010    1000001000011011    1000001000011100    1000001000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33305 - 33309

  --1000001000011110    1000001000011111    1000001000100000    1000001000100001    1000001000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33310 - 33314

  --1000001000100011    1000001000100100    1000001000100101    1000001000100110    1000001000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33315 - 33319

  --1000001000101000    1000001000101001    1000001000101010    1000001000101011    1000001000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33320 - 33324

  --1000001000101101    1000001000101110    1000001000101111    1000001000110000    1000001000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33325 - 33329

  --1000001000110010    1000001000110011    1000001000110100    1000001000110101    1000001000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33330 - 33334

  --1000001000110111    1000001000111000    1000001000111001    1000001000111010    1000001000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33335 - 33339

  --1000001000111100    1000001000111101    1000001000111110    1000001000111111    1000001001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33340 - 33344

  --1000001001000001    1000001001000010    1000001001000011    1000001001000100    1000001001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33345 - 33349

  --1000001001000110    1000001001000111    1000001001001000    1000001001001001    1000001001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33350 - 33354

  --1000001001001011    1000001001001100    1000001001001101    1000001001001110    1000001001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33355 - 33359

  --1000001001010000    1000001001010001    1000001001010010    1000001001010011    1000001001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33360 - 33364

  --1000001001010101    1000001001010110    1000001001010111    1000001001011000    1000001001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33365 - 33369

  --1000001001011010    1000001001011011    1000001001011100    1000001001011101    1000001001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33370 - 33374

  --1000001001011111    1000001001100000    1000001001100001    1000001001100010    1000001001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33375 - 33379

  --1000001001100100    1000001001100101    1000001001100110    1000001001100111    1000001001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33380 - 33384

  --1000001001101001    1000001001101010    1000001001101011    1000001001101100    1000001001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33385 - 33389

  --1000001001101110    1000001001101111    1000001001110000    1000001001110001    1000001001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33390 - 33394

  --1000001001110011    1000001001110100    1000001001110101    1000001001110110    1000001001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33395 - 33399

  --1000001001111000    1000001001111001    1000001001111010    1000001001111011    1000001001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33400 - 33404

  --1000001001111101    1000001001111110    1000001001111111    1000001010000000    1000001010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33405 - 33409

  --1000001010000010    1000001010000011    1000001010000100    1000001010000101    1000001010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33410 - 33414

  --1000001010000111    1000001010001000    1000001010001001    1000001010001010    1000001010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33415 - 33419

  --1000001010001100    1000001010001101    1000001010001110    1000001010001111    1000001010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33420 - 33424

  --1000001010010001    1000001010010010    1000001010010011    1000001010010100    1000001010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33425 - 33429

  --1000001010010110    1000001010010111    1000001010011000    1000001010011001    1000001010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33430 - 33434

  --1000001010011011    1000001010011100    1000001010011101    1000001010011110    1000001010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33435 - 33439

  --1000001010100000    1000001010100001    1000001010100010    1000001010100011    1000001010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33440 - 33444

  --1000001010100101    1000001010100110    1000001010100111    1000001010101000    1000001010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33445 - 33449

  --1000001010101010    1000001010101011    1000001010101100    1000001010101101    1000001010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33450 - 33454

  --1000001010101111    1000001010110000    1000001010110001    1000001010110010    1000001010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33455 - 33459

  --1000001010110100    1000001010110101    1000001010110110    1000001010110111    1000001010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33460 - 33464

  --1000001010111001    1000001010111010    1000001010111011    1000001010111100    1000001010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33465 - 33469

  --1000001010111110    1000001010111111    1000001011000000    1000001011000001    1000001011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33470 - 33474

  --1000001011000011    1000001011000100    1000001011000101    1000001011000110    1000001011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33475 - 33479

  --1000001011001000    1000001011001001    1000001011001010    1000001011001011    1000001011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33480 - 33484

  --1000001011001101    1000001011001110    1000001011001111    1000001011010000    1000001011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33485 - 33489

  --1000001011010010    1000001011010011    1000001011010100    1000001011010101    1000001011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33490 - 33494

  --1000001011010111    1000001011011000    1000001011011001    1000001011011010    1000001011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33495 - 33499

  --1000001011011100    1000001011011101    1000001011011110    1000001011011111    1000001011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33500 - 33504

  --1000001011100001    1000001011100010    1000001011100011    1000001011100100    1000001011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33505 - 33509

  --1000001011100110    1000001011100111    1000001011101000    1000001011101001    1000001011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33510 - 33514

  --1000001011101011    1000001011101100    1000001011101101    1000001011101110    1000001011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33515 - 33519

  --1000001011110000    1000001011110001    1000001011110010    1000001011110011    1000001011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33520 - 33524

  --1000001011110101    1000001011110110    1000001011110111    1000001011111000    1000001011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33525 - 33529

  --1000001011111010    1000001011111011    1000001011111100    1000001011111101    1000001011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33530 - 33534

  --1000001011111111    1000001100000000    1000001100000001    1000001100000010    1000001100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33535 - 33539

  --1000001100000100    1000001100000101    1000001100000110    1000001100000111    1000001100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33540 - 33544

  --1000001100001001    1000001100001010    1000001100001011    1000001100001100    1000001100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33545 - 33549

  --1000001100001110    1000001100001111    1000001100010000    1000001100010001    1000001100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33550 - 33554

  --1000001100010011    1000001100010100    1000001100010101    1000001100010110    1000001100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33555 - 33559

  --1000001100011000    1000001100011001    1000001100011010    1000001100011011    1000001100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33560 - 33564

  --1000001100011101    1000001100011110    1000001100011111    1000001100100000    1000001100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33565 - 33569

  --1000001100100010    1000001100100011    1000001100100100    1000001100100101    1000001100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33570 - 33574

  --1000001100100111    1000001100101000    1000001100101001    1000001100101010    1000001100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33575 - 33579

  --1000001100101100    1000001100101101    1000001100101110    1000001100101111    1000001100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33580 - 33584

  --1000001100110001    1000001100110010    1000001100110011    1000001100110100    1000001100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33585 - 33589

  --1000001100110110    1000001100110111    1000001100111000    1000001100111001    1000001100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33590 - 33594

  --1000001100111011    1000001100111100    1000001100111101    1000001100111110    1000001100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33595 - 33599

  --1000001101000000    1000001101000001    1000001101000010    1000001101000011    1000001101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33600 - 33604

  --1000001101000101    1000001101000110    1000001101000111    1000001101001000    1000001101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33605 - 33609

  --1000001101001010    1000001101001011    1000001101001100    1000001101001101    1000001101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33610 - 33614

  --1000001101001111    1000001101010000    1000001101010001    1000001101010010    1000001101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33615 - 33619

  --1000001101010100    1000001101010101    1000001101010110    1000001101010111    1000001101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33620 - 33624

  --1000001101011001    1000001101011010    1000001101011011    1000001101011100    1000001101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33625 - 33629

  --1000001101011110    1000001101011111    1000001101100000    1000001101100001    1000001101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33630 - 33634

  --1000001101100011    1000001101100100    1000001101100101    1000001101100110    1000001101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33635 - 33639

  --1000001101101000    1000001101101001    1000001101101010    1000001101101011    1000001101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33640 - 33644

  --1000001101101101    1000001101101110    1000001101101111    1000001101110000    1000001101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33645 - 33649

  --1000001101110010    1000001101110011    1000001101110100    1000001101110101    1000001101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33650 - 33654

  --1000001101110111    1000001101111000    1000001101111001    1000001101111010    1000001101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33655 - 33659

  --1000001101111100    1000001101111101    1000001101111110    1000001101111111    1000001110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33660 - 33664

  --1000001110000001    1000001110000010    1000001110000011    1000001110000100    1000001110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33665 - 33669

  --1000001110000110    1000001110000111    1000001110001000    1000001110001001    1000001110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33670 - 33674

  --1000001110001011    1000001110001100    1000001110001101    1000001110001110    1000001110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33675 - 33679

  --1000001110010000    1000001110010001    1000001110010010    1000001110010011    1000001110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33680 - 33684

  --1000001110010101    1000001110010110    1000001110010111    1000001110011000    1000001110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33685 - 33689

  --1000001110011010    1000001110011011    1000001110011100    1000001110011101    1000001110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33690 - 33694

  --1000001110011111    1000001110100000    1000001110100001    1000001110100010    1000001110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33695 - 33699

  --1000001110100100    1000001110100101    1000001110100110    1000001110100111    1000001110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33700 - 33704

  --1000001110101001    1000001110101010    1000001110101011    1000001110101100    1000001110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33705 - 33709

  --1000001110101110    1000001110101111    1000001110110000    1000001110110001    1000001110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33710 - 33714

  --1000001110110011    1000001110110100    1000001110110101    1000001110110110    1000001110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33715 - 33719

  --1000001110111000    1000001110111001    1000001110111010    1000001110111011    1000001110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33720 - 33724

  --1000001110111101    1000001110111110    1000001110111111    1000001111000000    1000001111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33725 - 33729

  --1000001111000010    1000001111000011    1000001111000100    1000001111000101    1000001111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33730 - 33734

  --1000001111000111    1000001111001000    1000001111001001    1000001111001010    1000001111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33735 - 33739

  --1000001111001100    1000001111001101    1000001111001110    1000001111001111    1000001111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33740 - 33744

  --1000001111010001    1000001111010010    1000001111010011    1000001111010100    1000001111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33745 - 33749

  --1000001111010110    1000001111010111    1000001111011000    1000001111011001    1000001111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33750 - 33754

  --1000001111011011    1000001111011100    1000001111011101    1000001111011110    1000001111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33755 - 33759

  --1000001111100000    1000001111100001    1000001111100010    1000001111100011    1000001111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33760 - 33764

  --1000001111100101    1000001111100110    1000001111100111    1000001111101000    1000001111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33765 - 33769

  --1000001111101010    1000001111101011    1000001111101100    1000001111101101    1000001111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33770 - 33774

  --1000001111101111    1000001111110000    1000001111110001    1000001111110010    1000001111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33775 - 33779

  --1000001111110100    1000001111110101    1000001111110110    1000001111110111    1000001111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33780 - 33784

  --1000001111111001    1000001111111010    1000001111111011    1000001111111100    1000001111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33785 - 33789

  --1000001111111110    1000001111111111    1000010000000000    1000010000000001    1000010000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33790 - 33794

  --1000010000000011    1000010000000100    1000010000000101    1000010000000110    1000010000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33795 - 33799

  --1000010000001000    1000010000001001    1000010000001010    1000010000001011    1000010000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33800 - 33804

  --1000010000001101    1000010000001110    1000010000001111    1000010000010000    1000010000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33805 - 33809

  --1000010000010010    1000010000010011    1000010000010100    1000010000010101    1000010000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33810 - 33814

  --1000010000010111    1000010000011000    1000010000011001    1000010000011010    1000010000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33815 - 33819

  --1000010000011100    1000010000011101    1000010000011110    1000010000011111    1000010000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33820 - 33824

  --1000010000100001    1000010000100010    1000010000100011    1000010000100100    1000010000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33825 - 33829

  --1000010000100110    1000010000100111    1000010000101000    1000010000101001    1000010000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33830 - 33834

  --1000010000101011    1000010000101100    1000010000101101    1000010000101110    1000010000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33835 - 33839

  --1000010000110000    1000010000110001    1000010000110010    1000010000110011    1000010000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33840 - 33844

  --1000010000110101    1000010000110110    1000010000110111    1000010000111000    1000010000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33845 - 33849

  --1000010000111010    1000010000111011    1000010000111100    1000010000111101    1000010000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33850 - 33854

  --1000010000111111    1000010001000000    1000010001000001    1000010001000010    1000010001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33855 - 33859

  --1000010001000100    1000010001000101    1000010001000110    1000010001000111    1000010001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33860 - 33864

  --1000010001001001    1000010001001010    1000010001001011    1000010001001100    1000010001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33865 - 33869

  --1000010001001110    1000010001001111    1000010001010000    1000010001010001    1000010001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33870 - 33874

  --1000010001010011    1000010001010100    1000010001010101    1000010001010110    1000010001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33875 - 33879

  --1000010001011000    1000010001011001    1000010001011010    1000010001011011    1000010001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33880 - 33884

  --1000010001011101    1000010001011110    1000010001011111    1000010001100000    1000010001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33885 - 33889

  --1000010001100010    1000010001100011    1000010001100100    1000010001100101    1000010001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33890 - 33894

  --1000010001100111    1000010001101000    1000010001101001    1000010001101010    1000010001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33895 - 33899

  --1000010001101100    1000010001101101    1000010001101110    1000010001101111    1000010001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33900 - 33904

  --1000010001110001    1000010001110010    1000010001110011    1000010001110100    1000010001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33905 - 33909

  --1000010001110110    1000010001110111    1000010001111000    1000010001111001    1000010001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33910 - 33914

  --1000010001111011    1000010001111100    1000010001111101    1000010001111110    1000010001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33915 - 33919

  --1000010010000000    1000010010000001    1000010010000010    1000010010000011    1000010010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33920 - 33924

  --1000010010000101    1000010010000110    1000010010000111    1000010010001000    1000010010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33925 - 33929

  --1000010010001010    1000010010001011    1000010010001100    1000010010001101    1000010010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33930 - 33934

  --1000010010001111    1000010010010000    1000010010010001    1000010010010010    1000010010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33935 - 33939

  --1000010010010100    1000010010010101    1000010010010110    1000010010010111    1000010010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33940 - 33944

  --1000010010011001    1000010010011010    1000010010011011    1000010010011100    1000010010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33945 - 33949

  --1000010010011110    1000010010011111    1000010010100000    1000010010100001    1000010010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33950 - 33954

  --1000010010100011    1000010010100100    1000010010100101    1000010010100110    1000010010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33955 - 33959

  --1000010010101000    1000010010101001    1000010010101010    1000010010101011    1000010010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33960 - 33964

  --1000010010101101    1000010010101110    1000010010101111    1000010010110000    1000010010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33965 - 33969

  --1000010010110010    1000010010110011    1000010010110100    1000010010110101    1000010010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33970 - 33974

  --1000010010110111    1000010010111000    1000010010111001    1000010010111010    1000010010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33975 - 33979

  --1000010010111100    1000010010111101    1000010010111110    1000010010111111    1000010011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33980 - 33984

  --1000010011000001    1000010011000010    1000010011000011    1000010011000100    1000010011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33985 - 33989

  --1000010011000110    1000010011000111    1000010011001000    1000010011001001    1000010011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33990 - 33994

  --1000010011001011    1000010011001100    1000010011001101    1000010011001110    1000010011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 33995 - 33999

  --1000010011010000    1000010011010001    1000010011010010    1000010011010011    1000010011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34000 - 34004

  --1000010011010101    1000010011010110    1000010011010111    1000010011011000    1000010011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34005 - 34009

  --1000010011011010    1000010011011011    1000010011011100    1000010011011101    1000010011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34010 - 34014

  --1000010011011111    1000010011100000    1000010011100001    1000010011100010    1000010011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34015 - 34019

  --1000010011100100    1000010011100101    1000010011100110    1000010011100111    1000010011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34020 - 34024

  --1000010011101001    1000010011101010    1000010011101011    1000010011101100    1000010011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34025 - 34029

  --1000010011101110    1000010011101111    1000010011110000    1000010011110001    1000010011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34030 - 34034

  --1000010011110011    1000010011110100    1000010011110101    1000010011110110    1000010011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34035 - 34039

  --1000010011111000    1000010011111001    1000010011111010    1000010011111011    1000010011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34040 - 34044

  --1000010011111101    1000010011111110    1000010011111111    1000010100000000    1000010100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34045 - 34049

  --1000010100000010    1000010100000011    1000010100000100    1000010100000101    1000010100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34050 - 34054

  --1000010100000111    1000010100001000    1000010100001001    1000010100001010    1000010100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34055 - 34059

  --1000010100001100    1000010100001101    1000010100001110    1000010100001111    1000010100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34060 - 34064

  --1000010100010001    1000010100010010    1000010100010011    1000010100010100    1000010100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34065 - 34069

  --1000010100010110    1000010100010111    1000010100011000    1000010100011001    1000010100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34070 - 34074

  --1000010100011011    1000010100011100    1000010100011101    1000010100011110    1000010100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34075 - 34079

  --1000010100100000    1000010100100001    1000010100100010    1000010100100011    1000010100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34080 - 34084

  --1000010100100101    1000010100100110    1000010100100111    1000010100101000    1000010100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34085 - 34089

  --1000010100101010    1000010100101011    1000010100101100    1000010100101101    1000010100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34090 - 34094

  --1000010100101111    1000010100110000    1000010100110001    1000010100110010    1000010100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34095 - 34099

  --1000010100110100    1000010100110101    1000010100110110    1000010100110111    1000010100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34100 - 34104

  --1000010100111001    1000010100111010    1000010100111011    1000010100111100    1000010100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34105 - 34109

  --1000010100111110    1000010100111111    1000010101000000    1000010101000001    1000010101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34110 - 34114

  --1000010101000011    1000010101000100    1000010101000101    1000010101000110    1000010101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34115 - 34119

  --1000010101001000    1000010101001001    1000010101001010    1000010101001011    1000010101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34120 - 34124

  --1000010101001101    1000010101001110    1000010101001111    1000010101010000    1000010101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34125 - 34129

  --1000010101010010    1000010101010011    1000010101010100    1000010101010101    1000010101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34130 - 34134

  --1000010101010111    1000010101011000    1000010101011001    1000010101011010    1000010101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34135 - 34139

  --1000010101011100    1000010101011101    1000010101011110    1000010101011111    1000010101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34140 - 34144

  --1000010101100001    1000010101100010    1000010101100011    1000010101100100    1000010101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34145 - 34149

  --1000010101100110    1000010101100111    1000010101101000    1000010101101001    1000010101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34150 - 34154

  --1000010101101011    1000010101101100    1000010101101101    1000010101101110    1000010101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34155 - 34159

  --1000010101110000    1000010101110001    1000010101110010    1000010101110011    1000010101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34160 - 34164

  --1000010101110101    1000010101110110    1000010101110111    1000010101111000    1000010101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34165 - 34169

  --1000010101111010    1000010101111011    1000010101111100    1000010101111101    1000010101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34170 - 34174

  --1000010101111111    1000010110000000    1000010110000001    1000010110000010    1000010110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34175 - 34179

  --1000010110000100    1000010110000101    1000010110000110    1000010110000111    1000010110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34180 - 34184

  --1000010110001001    1000010110001010    1000010110001011    1000010110001100    1000010110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34185 - 34189

  --1000010110001110    1000010110001111    1000010110010000    1000010110010001    1000010110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34190 - 34194

  --1000010110010011    1000010110010100    1000010110010101    1000010110010110    1000010110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34195 - 34199

  --1000010110011000    1000010110011001    1000010110011010    1000010110011011    1000010110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34200 - 34204

  --1000010110011101    1000010110011110    1000010110011111    1000010110100000    1000010110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34205 - 34209

  --1000010110100010    1000010110100011    1000010110100100    1000010110100101    1000010110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34210 - 34214

  --1000010110100111    1000010110101000    1000010110101001    1000010110101010    1000010110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34215 - 34219

  --1000010110101100    1000010110101101    1000010110101110    1000010110101111    1000010110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34220 - 34224

  --1000010110110001    1000010110110010    1000010110110011    1000010110110100    1000010110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34225 - 34229

  --1000010110110110    1000010110110111    1000010110111000    1000010110111001    1000010110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34230 - 34234

  --1000010110111011    1000010110111100    1000010110111101    1000010110111110    1000010110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34235 - 34239

  --1000010111000000    1000010111000001    1000010111000010    1000010111000011    1000010111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34240 - 34244

  --1000010111000101    1000010111000110    1000010111000111    1000010111001000    1000010111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34245 - 34249

  --1000010111001010    1000010111001011    1000010111001100    1000010111001101    1000010111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34250 - 34254

  --1000010111001111    1000010111010000    1000010111010001    1000010111010010    1000010111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34255 - 34259

  --1000010111010100    1000010111010101    1000010111010110    1000010111010111    1000010111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34260 - 34264

  --1000010111011001    1000010111011010    1000010111011011    1000010111011100    1000010111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34265 - 34269

  --1000010111011110    1000010111011111    1000010111100000    1000010111100001    1000010111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34270 - 34274

  --1000010111100011    1000010111100100    1000010111100101    1000010111100110    1000010111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34275 - 34279

  --1000010111101000    1000010111101001    1000010111101010    1000010111101011    1000010111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34280 - 34284

  --1000010111101101    1000010111101110    1000010111101111    1000010111110000    1000010111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34285 - 34289

  --1000010111110010    1000010111110011    1000010111110100    1000010111110101    1000010111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34290 - 34294

  --1000010111110111    1000010111111000    1000010111111001    1000010111111010    1000010111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34295 - 34299

  --1000010111111100    1000010111111101    1000010111111110    1000010111111111    1000011000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34300 - 34304

  --1000011000000001    1000011000000010    1000011000000011    1000011000000100    1000011000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34305 - 34309

  --1000011000000110    1000011000000111    1000011000001000    1000011000001001    1000011000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34310 - 34314

  --1000011000001011    1000011000001100    1000011000001101    1000011000001110    1000011000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34315 - 34319

  --1000011000010000    1000011000010001    1000011000010010    1000011000010011    1000011000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34320 - 34324

  --1000011000010101    1000011000010110    1000011000010111    1000011000011000    1000011000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34325 - 34329

  --1000011000011010    1000011000011011    1000011000011100    1000011000011101    1000011000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34330 - 34334

  --1000011000011111    1000011000100000    1000011000100001    1000011000100010    1000011000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34335 - 34339

  --1000011000100100    1000011000100101    1000011000100110    1000011000100111    1000011000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34340 - 34344

  --1000011000101001    1000011000101010    1000011000101011    1000011000101100    1000011000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34345 - 34349

  --1000011000101110    1000011000101111    1000011000110000    1000011000110001    1000011000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34350 - 34354

  --1000011000110011    1000011000110100    1000011000110101    1000011000110110    1000011000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34355 - 34359

  --1000011000111000    1000011000111001    1000011000111010    1000011000111011    1000011000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34360 - 34364

  --1000011000111101    1000011000111110    1000011000111111    1000011001000000    1000011001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34365 - 34369

  --1000011001000010    1000011001000011    1000011001000100    1000011001000101    1000011001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34370 - 34374

  --1000011001000111    1000011001001000    1000011001001001    1000011001001010    1000011001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34375 - 34379

  --1000011001001100    1000011001001101    1000011001001110    1000011001001111    1000011001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34380 - 34384

  --1000011001010001    1000011001010010    1000011001010011    1000011001010100    1000011001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34385 - 34389

  --1000011001010110    1000011001010111    1000011001011000    1000011001011001    1000011001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34390 - 34394

  --1000011001011011    1000011001011100    1000011001011101    1000011001011110    1000011001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34395 - 34399

  --1000011001100000    1000011001100001    1000011001100010    1000011001100011    1000011001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34400 - 34404

  --1000011001100101    1000011001100110    1000011001100111    1000011001101000    1000011001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34405 - 34409

  --1000011001101010    1000011001101011    1000011001101100    1000011001101101    1000011001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34410 - 34414

  --1000011001101111    1000011001110000    1000011001110001    1000011001110010    1000011001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34415 - 34419

  --1000011001110100    1000011001110101    1000011001110110    1000011001110111    1000011001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34420 - 34424

  --1000011001111001    1000011001111010    1000011001111011    1000011001111100    1000011001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34425 - 34429

  --1000011001111110    1000011001111111    1000011010000000    1000011010000001    1000011010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34430 - 34434

  --1000011010000011    1000011010000100    1000011010000101    1000011010000110    1000011010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34435 - 34439

  --1000011010001000    1000011010001001    1000011010001010    1000011010001011    1000011010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34440 - 34444

  --1000011010001101    1000011010001110    1000011010001111    1000011010010000    1000011010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34445 - 34449

  --1000011010010010    1000011010010011    1000011010010100    1000011010010101    1000011010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34450 - 34454

  --1000011010010111    1000011010011000    1000011010011001    1000011010011010    1000011010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34455 - 34459

  --1000011010011100    1000011010011101    1000011010011110    1000011010011111    1000011010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34460 - 34464

  --1000011010100001    1000011010100010    1000011010100011    1000011010100100    1000011010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34465 - 34469

  --1000011010100110    1000011010100111    1000011010101000    1000011010101001    1000011010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34470 - 34474

  --1000011010101011    1000011010101100    1000011010101101    1000011010101110    1000011010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34475 - 34479

  --1000011010110000    1000011010110001    1000011010110010    1000011010110011    1000011010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34480 - 34484

  --1000011010110101    1000011010110110    1000011010110111    1000011010111000    1000011010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34485 - 34489

  --1000011010111010    1000011010111011    1000011010111100    1000011010111101    1000011010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34490 - 34494

  --1000011010111111    1000011011000000    1000011011000001    1000011011000010    1000011011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34495 - 34499

  --1000011011000100    1000011011000101    1000011011000110    1000011011000111    1000011011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34500 - 34504

  --1000011011001001    1000011011001010    1000011011001011    1000011011001100    1000011011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34505 - 34509

  --1000011011001110    1000011011001111    1000011011010000    1000011011010001    1000011011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34510 - 34514

  --1000011011010011    1000011011010100    1000011011010101    1000011011010110    1000011011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34515 - 34519

  --1000011011011000    1000011011011001    1000011011011010    1000011011011011    1000011011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34520 - 34524

  --1000011011011101    1000011011011110    1000011011011111    1000011011100000    1000011011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34525 - 34529

  --1000011011100010    1000011011100011    1000011011100100    1000011011100101    1000011011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34530 - 34534

  --1000011011100111    1000011011101000    1000011011101001    1000011011101010    1000011011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34535 - 34539

  --1000011011101100    1000011011101101    1000011011101110    1000011011101111    1000011011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34540 - 34544

  --1000011011110001    1000011011110010    1000011011110011    1000011011110100    1000011011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34545 - 34549

  --1000011011110110    1000011011110111    1000011011111000    1000011011111001    1000011011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34550 - 34554

  --1000011011111011    1000011011111100    1000011011111101    1000011011111110    1000011011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34555 - 34559

  --1000011100000000    1000011100000001    1000011100000010    1000011100000011    1000011100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34560 - 34564

  --1000011100000101    1000011100000110    1000011100000111    1000011100001000    1000011100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34565 - 34569

  --1000011100001010    1000011100001011    1000011100001100    1000011100001101    1000011100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34570 - 34574

  --1000011100001111    1000011100010000    1000011100010001    1000011100010010    1000011100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34575 - 34579

  --1000011100010100    1000011100010101    1000011100010110    1000011100010111    1000011100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34580 - 34584

  --1000011100011001    1000011100011010    1000011100011011    1000011100011100    1000011100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34585 - 34589

  --1000011100011110    1000011100011111    1000011100100000    1000011100100001    1000011100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34590 - 34594

  --1000011100100011    1000011100100100    1000011100100101    1000011100100110    1000011100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34595 - 34599

  --1000011100101000    1000011100101001    1000011100101010    1000011100101011    1000011100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34600 - 34604

  --1000011100101101    1000011100101110    1000011100101111    1000011100110000    1000011100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34605 - 34609

  --1000011100110010    1000011100110011    1000011100110100    1000011100110101    1000011100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34610 - 34614

  --1000011100110111    1000011100111000    1000011100111001    1000011100111010    1000011100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34615 - 34619

  --1000011100111100    1000011100111101    1000011100111110    1000011100111111    1000011101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34620 - 34624

  --1000011101000001    1000011101000010    1000011101000011    1000011101000100    1000011101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34625 - 34629

  --1000011101000110    1000011101000111    1000011101001000    1000011101001001    1000011101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34630 - 34634

  --1000011101001011    1000011101001100    1000011101001101    1000011101001110    1000011101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34635 - 34639

  --1000011101010000    1000011101010001    1000011101010010    1000011101010011    1000011101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34640 - 34644

  --1000011101010101    1000011101010110    1000011101010111    1000011101011000    1000011101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34645 - 34649

  --1000011101011010    1000011101011011    1000011101011100    1000011101011101    1000011101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34650 - 34654

  --1000011101011111    1000011101100000    1000011101100001    1000011101100010    1000011101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34655 - 34659

  --1000011101100100    1000011101100101    1000011101100110    1000011101100111    1000011101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34660 - 34664

  --1000011101101001    1000011101101010    1000011101101011    1000011101101100    1000011101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34665 - 34669

  --1000011101101110    1000011101101111    1000011101110000    1000011101110001    1000011101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34670 - 34674

  --1000011101110011    1000011101110100    1000011101110101    1000011101110110    1000011101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34675 - 34679

  --1000011101111000    1000011101111001    1000011101111010    1000011101111011    1000011101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34680 - 34684

  --1000011101111101    1000011101111110    1000011101111111    1000011110000000    1000011110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34685 - 34689

  --1000011110000010    1000011110000011    1000011110000100    1000011110000101    1000011110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34690 - 34694

  --1000011110000111    1000011110001000    1000011110001001    1000011110001010    1000011110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34695 - 34699

  --1000011110001100    1000011110001101    1000011110001110    1000011110001111    1000011110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34700 - 34704

  --1000011110010001    1000011110010010    1000011110010011    1000011110010100    1000011110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34705 - 34709

  --1000011110010110    1000011110010111    1000011110011000    1000011110011001    1000011110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34710 - 34714

  --1000011110011011    1000011110011100    1000011110011101    1000011110011110    1000011110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34715 - 34719

  --1000011110100000    1000011110100001    1000011110100010    1000011110100011    1000011110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34720 - 34724

  --1000011110100101    1000011110100110    1000011110100111    1000011110101000    1000011110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34725 - 34729

  --1000011110101010    1000011110101011    1000011110101100    1000011110101101    1000011110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34730 - 34734

  --1000011110101111    1000011110110000    1000011110110001    1000011110110010    1000011110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34735 - 34739

  --1000011110110100    1000011110110101    1000011110110110    1000011110110111    1000011110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34740 - 34744

  --1000011110111001    1000011110111010    1000011110111011    1000011110111100    1000011110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34745 - 34749

  --1000011110111110    1000011110111111    1000011111000000    1000011111000001    1000011111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34750 - 34754

  --1000011111000011    1000011111000100    1000011111000101    1000011111000110    1000011111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34755 - 34759

  --1000011111001000    1000011111001001    1000011111001010    1000011111001011    1000011111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34760 - 34764

  --1000011111001101    1000011111001110    1000011111001111    1000011111010000    1000011111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34765 - 34769

  --1000011111010010    1000011111010011    1000011111010100    1000011111010101    1000011111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34770 - 34774

  --1000011111010111    1000011111011000    1000011111011001    1000011111011010    1000011111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34775 - 34779

  --1000011111011100    1000011111011101    1000011111011110    1000011111011111    1000011111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34780 - 34784

  --1000011111100001    1000011111100010    1000011111100011    1000011111100100    1000011111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34785 - 34789

  --1000011111100110    1000011111100111    1000011111101000    1000011111101001    1000011111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34790 - 34794

  --1000011111101011    1000011111101100    1000011111101101    1000011111101110    1000011111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34795 - 34799

  --1000011111110000    1000011111110001    1000011111110010    1000011111110011    1000011111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34800 - 34804

  --1000011111110101    1000011111110110    1000011111110111    1000011111111000    1000011111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34805 - 34809

  --1000011111111010    1000011111111011    1000011111111100    1000011111111101    1000011111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34810 - 34814

  --1000011111111111    1000100000000000    1000100000000001    1000100000000010    1000100000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34815 - 34819

  --1000100000000100    1000100000000101    1000100000000110    1000100000000111    1000100000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34820 - 34824

  --1000100000001001    1000100000001010    1000100000001011    1000100000001100    1000100000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34825 - 34829

  --1000100000001110    1000100000001111    1000100000010000    1000100000010001    1000100000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34830 - 34834

  --1000100000010011    1000100000010100    1000100000010101    1000100000010110    1000100000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34835 - 34839

  --1000100000011000    1000100000011001    1000100000011010    1000100000011011    1000100000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34840 - 34844

  --1000100000011101    1000100000011110    1000100000011111    1000100000100000    1000100000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34845 - 34849

  --1000100000100010    1000100000100011    1000100000100100    1000100000100101    1000100000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34850 - 34854

  --1000100000100111    1000100000101000    1000100000101001    1000100000101010    1000100000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34855 - 34859

  --1000100000101100    1000100000101101    1000100000101110    1000100000101111    1000100000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34860 - 34864

  --1000100000110001    1000100000110010    1000100000110011    1000100000110100    1000100000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34865 - 34869

  --1000100000110110    1000100000110111    1000100000111000    1000100000111001    1000100000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34870 - 34874

  --1000100000111011    1000100000111100    1000100000111101    1000100000111110    1000100000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34875 - 34879

  --1000100001000000    1000100001000001    1000100001000010    1000100001000011    1000100001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34880 - 34884

  --1000100001000101    1000100001000110    1000100001000111    1000100001001000    1000100001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34885 - 34889

  --1000100001001010    1000100001001011    1000100001001100    1000100001001101    1000100001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34890 - 34894

  --1000100001001111    1000100001010000    1000100001010001    1000100001010010    1000100001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34895 - 34899

  --1000100001010100    1000100001010101    1000100001010110    1000100001010111    1000100001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34900 - 34904

  --1000100001011001    1000100001011010    1000100001011011    1000100001011100    1000100001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34905 - 34909

  --1000100001011110    1000100001011111    1000100001100000    1000100001100001    1000100001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34910 - 34914

  --1000100001100011    1000100001100100    1000100001100101    1000100001100110    1000100001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34915 - 34919

  --1000100001101000    1000100001101001    1000100001101010    1000100001101011    1000100001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34920 - 34924

  --1000100001101101    1000100001101110    1000100001101111    1000100001110000    1000100001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34925 - 34929

  --1000100001110010    1000100001110011    1000100001110100    1000100001110101    1000100001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34930 - 34934

  --1000100001110111    1000100001111000    1000100001111001    1000100001111010    1000100001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34935 - 34939

  --1000100001111100    1000100001111101    1000100001111110    1000100001111111    1000100010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34940 - 34944

  --1000100010000001    1000100010000010    1000100010000011    1000100010000100    1000100010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34945 - 34949

  --1000100010000110    1000100010000111    1000100010001000    1000100010001001    1000100010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34950 - 34954

  --1000100010001011    1000100010001100    1000100010001101    1000100010001110    1000100010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34955 - 34959

  --1000100010010000    1000100010010001    1000100010010010    1000100010010011    1000100010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34960 - 34964

  --1000100010010101    1000100010010110    1000100010010111    1000100010011000    1000100010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34965 - 34969

  --1000100010011010    1000100010011011    1000100010011100    1000100010011101    1000100010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34970 - 34974

  --1000100010011111    1000100010100000    1000100010100001    1000100010100010    1000100010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34975 - 34979

  --1000100010100100    1000100010100101    1000100010100110    1000100010100111    1000100010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34980 - 34984

  --1000100010101001    1000100010101010    1000100010101011    1000100010101100    1000100010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34985 - 34989

  --1000100010101110    1000100010101111    1000100010110000    1000100010110001    1000100010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34990 - 34994

  --1000100010110011    1000100010110100    1000100010110101    1000100010110110    1000100010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 34995 - 34999

  --1000100010111000    1000100010111001    1000100010111010    1000100010111011    1000100010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35000 - 35004

  --1000100010111101    1000100010111110    1000100010111111    1000100011000000    1000100011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35005 - 35009

  --1000100011000010    1000100011000011    1000100011000100    1000100011000101    1000100011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35010 - 35014

  --1000100011000111    1000100011001000    1000100011001001    1000100011001010    1000100011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35015 - 35019

  --1000100011001100    1000100011001101    1000100011001110    1000100011001111    1000100011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35020 - 35024

  --1000100011010001    1000100011010010    1000100011010011    1000100011010100    1000100011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35025 - 35029

  --1000100011010110    1000100011010111    1000100011011000    1000100011011001    1000100011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35030 - 35034

  --1000100011011011    1000100011011100    1000100011011101    1000100011011110    1000100011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35035 - 35039

  --1000100011100000    1000100011100001    1000100011100010    1000100011100011    1000100011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35040 - 35044

  --1000100011100101    1000100011100110    1000100011100111    1000100011101000    1000100011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35045 - 35049

  --1000100011101010    1000100011101011    1000100011101100    1000100011101101    1000100011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35050 - 35054

  --1000100011101111    1000100011110000    1000100011110001    1000100011110010    1000100011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35055 - 35059

  --1000100011110100    1000100011110101    1000100011110110    1000100011110111    1000100011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35060 - 35064

  --1000100011111001    1000100011111010    1000100011111011    1000100011111100    1000100011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35065 - 35069

  --1000100011111110    1000100011111111    1000100100000000    1000100100000001    1000100100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35070 - 35074

  --1000100100000011    1000100100000100    1000100100000101    1000100100000110    1000100100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35075 - 35079

  --1000100100001000    1000100100001001    1000100100001010    1000100100001011    1000100100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35080 - 35084

  --1000100100001101    1000100100001110    1000100100001111    1000100100010000    1000100100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35085 - 35089

  --1000100100010010    1000100100010011    1000100100010100    1000100100010101    1000100100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35090 - 35094

  --1000100100010111    1000100100011000    1000100100011001    1000100100011010    1000100100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35095 - 35099

  --1000100100011100    1000100100011101    1000100100011110    1000100100011111    1000100100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35100 - 35104

  --1000100100100001    1000100100100010    1000100100100011    1000100100100100    1000100100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35105 - 35109

  --1000100100100110    1000100100100111    1000100100101000    1000100100101001    1000100100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35110 - 35114

  --1000100100101011    1000100100101100    1000100100101101    1000100100101110    1000100100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35115 - 35119

  --1000100100110000    1000100100110001    1000100100110010    1000100100110011    1000100100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35120 - 35124

  --1000100100110101    1000100100110110    1000100100110111    1000100100111000    1000100100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35125 - 35129

  --1000100100111010    1000100100111011    1000100100111100    1000100100111101    1000100100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35130 - 35134

  --1000100100111111    1000100101000000    1000100101000001    1000100101000010    1000100101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35135 - 35139

  --1000100101000100    1000100101000101    1000100101000110    1000100101000111    1000100101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35140 - 35144

  --1000100101001001    1000100101001010    1000100101001011    1000100101001100    1000100101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35145 - 35149

  --1000100101001110    1000100101001111    1000100101010000    1000100101010001    1000100101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35150 - 35154

  --1000100101010011    1000100101010100    1000100101010101    1000100101010110    1000100101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35155 - 35159

  --1000100101011000    1000100101011001    1000100101011010    1000100101011011    1000100101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35160 - 35164

  --1000100101011101    1000100101011110    1000100101011111    1000100101100000    1000100101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35165 - 35169

  --1000100101100010    1000100101100011    1000100101100100    1000100101100101    1000100101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35170 - 35174

  --1000100101100111    1000100101101000    1000100101101001    1000100101101010    1000100101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35175 - 35179

  --1000100101101100    1000100101101101    1000100101101110    1000100101101111    1000100101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35180 - 35184

  --1000100101110001    1000100101110010    1000100101110011    1000100101110100    1000100101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35185 - 35189

  --1000100101110110    1000100101110111    1000100101111000    1000100101111001    1000100101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35190 - 35194

  --1000100101111011    1000100101111100    1000100101111101    1000100101111110    1000100101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35195 - 35199

  --1000100110000000    1000100110000001    1000100110000010    1000100110000011    1000100110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35200 - 35204

  --1000100110000101    1000100110000110    1000100110000111    1000100110001000    1000100110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35205 - 35209

  --1000100110001010    1000100110001011    1000100110001100    1000100110001101    1000100110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35210 - 35214

  --1000100110001111    1000100110010000    1000100110010001    1000100110010010    1000100110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35215 - 35219

  --1000100110010100    1000100110010101    1000100110010110    1000100110010111    1000100110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35220 - 35224

  --1000100110011001    1000100110011010    1000100110011011    1000100110011100    1000100110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35225 - 35229

  --1000100110011110    1000100110011111    1000100110100000    1000100110100001    1000100110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35230 - 35234

  --1000100110100011    1000100110100100    1000100110100101    1000100110100110    1000100110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35235 - 35239

  --1000100110101000    1000100110101001    1000100110101010    1000100110101011    1000100110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35240 - 35244

  --1000100110101101    1000100110101110    1000100110101111    1000100110110000    1000100110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35245 - 35249

  --1000100110110010    1000100110110011    1000100110110100    1000100110110101    1000100110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35250 - 35254

  --1000100110110111    1000100110111000    1000100110111001    1000100110111010    1000100110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35255 - 35259

  --1000100110111100    1000100110111101    1000100110111110    1000100110111111    1000100111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35260 - 35264

  --1000100111000001    1000100111000010    1000100111000011    1000100111000100    1000100111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35265 - 35269

  --1000100111000110    1000100111000111    1000100111001000    1000100111001001    1000100111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35270 - 35274

  --1000100111001011    1000100111001100    1000100111001101    1000100111001110    1000100111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35275 - 35279

  --1000100111010000    1000100111010001    1000100111010010    1000100111010011    1000100111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35280 - 35284

  --1000100111010101    1000100111010110    1000100111010111    1000100111011000    1000100111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35285 - 35289

  --1000100111011010    1000100111011011    1000100111011100    1000100111011101    1000100111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35290 - 35294

  --1000100111011111    1000100111100000    1000100111100001    1000100111100010    1000100111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35295 - 35299

  --1000100111100100    1000100111100101    1000100111100110    1000100111100111    1000100111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35300 - 35304

  --1000100111101001    1000100111101010    1000100111101011    1000100111101100    1000100111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35305 - 35309

  --1000100111101110    1000100111101111    1000100111110000    1000100111110001    1000100111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35310 - 35314

  --1000100111110011    1000100111110100    1000100111110101    1000100111110110    1000100111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35315 - 35319

  --1000100111111000    1000100111111001    1000100111111010    1000100111111011    1000100111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35320 - 35324

  --1000100111111101    1000100111111110    1000100111111111    1000101000000000    1000101000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35325 - 35329

  --1000101000000010    1000101000000011    1000101000000100    1000101000000101    1000101000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35330 - 35334

  --1000101000000111    1000101000001000    1000101000001001    1000101000001010    1000101000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35335 - 35339

  --1000101000001100    1000101000001101    1000101000001110    1000101000001111    1000101000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35340 - 35344

  --1000101000010001    1000101000010010    1000101000010011    1000101000010100    1000101000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35345 - 35349

  --1000101000010110    1000101000010111    1000101000011000    1000101000011001    1000101000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35350 - 35354

  --1000101000011011    1000101000011100    1000101000011101    1000101000011110    1000101000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35355 - 35359

  --1000101000100000    1000101000100001    1000101000100010    1000101000100011    1000101000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35360 - 35364

  --1000101000100101    1000101000100110    1000101000100111    1000101000101000    1000101000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35365 - 35369

  --1000101000101010    1000101000101011    1000101000101100    1000101000101101    1000101000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35370 - 35374

  --1000101000101111    1000101000110000    1000101000110001    1000101000110010    1000101000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35375 - 35379

  --1000101000110100    1000101000110101    1000101000110110    1000101000110111    1000101000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35380 - 35384

  --1000101000111001    1000101000111010    1000101000111011    1000101000111100    1000101000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35385 - 35389

  --1000101000111110    1000101000111111    1000101001000000    1000101001000001    1000101001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35390 - 35394

  --1000101001000011    1000101001000100    1000101001000101    1000101001000110    1000101001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35395 - 35399

  --1000101001001000    1000101001001001    1000101001001010    1000101001001011    1000101001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35400 - 35404

  --1000101001001101    1000101001001110    1000101001001111    1000101001010000    1000101001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35405 - 35409

  --1000101001010010    1000101001010011    1000101001010100    1000101001010101    1000101001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35410 - 35414

  --1000101001010111    1000101001011000    1000101001011001    1000101001011010    1000101001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35415 - 35419

  --1000101001011100    1000101001011101    1000101001011110    1000101001011111    1000101001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35420 - 35424

  --1000101001100001    1000101001100010    1000101001100011    1000101001100100    1000101001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35425 - 35429

  --1000101001100110    1000101001100111    1000101001101000    1000101001101001    1000101001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35430 - 35434

  --1000101001101011    1000101001101100    1000101001101101    1000101001101110    1000101001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35435 - 35439

  --1000101001110000    1000101001110001    1000101001110010    1000101001110011    1000101001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35440 - 35444

  --1000101001110101    1000101001110110    1000101001110111    1000101001111000    1000101001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35445 - 35449

  --1000101001111010    1000101001111011    1000101001111100    1000101001111101    1000101001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35450 - 35454

  --1000101001111111    1000101010000000    1000101010000001    1000101010000010    1000101010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35455 - 35459

  --1000101010000100    1000101010000101    1000101010000110    1000101010000111    1000101010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35460 - 35464

  --1000101010001001    1000101010001010    1000101010001011    1000101010001100    1000101010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35465 - 35469

  --1000101010001110    1000101010001111    1000101010010000    1000101010010001    1000101010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35470 - 35474

  --1000101010010011    1000101010010100    1000101010010101    1000101010010110    1000101010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35475 - 35479

  --1000101010011000    1000101010011001    1000101010011010    1000101010011011    1000101010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35480 - 35484

  --1000101010011101    1000101010011110    1000101010011111    1000101010100000    1000101010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35485 - 35489

  --1000101010100010    1000101010100011    1000101010100100    1000101010100101    1000101010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35490 - 35494

  --1000101010100111    1000101010101000    1000101010101001    1000101010101010    1000101010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35495 - 35499

  --1000101010101100    1000101010101101    1000101010101110    1000101010101111    1000101010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35500 - 35504

  --1000101010110001    1000101010110010    1000101010110011    1000101010110100    1000101010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35505 - 35509

  --1000101010110110    1000101010110111    1000101010111000    1000101010111001    1000101010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35510 - 35514

  --1000101010111011    1000101010111100    1000101010111101    1000101010111110    1000101010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35515 - 35519

  --1000101011000000    1000101011000001    1000101011000010    1000101011000011    1000101011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35520 - 35524

  --1000101011000101    1000101011000110    1000101011000111    1000101011001000    1000101011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35525 - 35529

  --1000101011001010    1000101011001011    1000101011001100    1000101011001101    1000101011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35530 - 35534

  --1000101011001111    1000101011010000    1000101011010001    1000101011010010    1000101011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35535 - 35539

  --1000101011010100    1000101011010101    1000101011010110    1000101011010111    1000101011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35540 - 35544

  --1000101011011001    1000101011011010    1000101011011011    1000101011011100    1000101011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35545 - 35549

  --1000101011011110    1000101011011111    1000101011100000    1000101011100001    1000101011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35550 - 35554

  --1000101011100011    1000101011100100    1000101011100101    1000101011100110    1000101011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35555 - 35559

  --1000101011101000    1000101011101001    1000101011101010    1000101011101011    1000101011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35560 - 35564

  --1000101011101101    1000101011101110    1000101011101111    1000101011110000    1000101011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35565 - 35569

  --1000101011110010    1000101011110011    1000101011110100    1000101011110101    1000101011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35570 - 35574

  --1000101011110111    1000101011111000    1000101011111001    1000101011111010    1000101011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35575 - 35579

  --1000101011111100    1000101011111101    1000101011111110    1000101011111111    1000101100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35580 - 35584

  --1000101100000001    1000101100000010    1000101100000011    1000101100000100    1000101100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35585 - 35589

  --1000101100000110    1000101100000111    1000101100001000    1000101100001001    1000101100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35590 - 35594

  --1000101100001011    1000101100001100    1000101100001101    1000101100001110    1000101100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35595 - 35599

  --1000101100010000    1000101100010001    1000101100010010    1000101100010011    1000101100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35600 - 35604

  --1000101100010101    1000101100010110    1000101100010111    1000101100011000    1000101100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35605 - 35609

  --1000101100011010    1000101100011011    1000101100011100    1000101100011101    1000101100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35610 - 35614

  --1000101100011111    1000101100100000    1000101100100001    1000101100100010    1000101100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35615 - 35619

  --1000101100100100    1000101100100101    1000101100100110    1000101100100111    1000101100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35620 - 35624

  --1000101100101001    1000101100101010    1000101100101011    1000101100101100    1000101100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35625 - 35629

  --1000101100101110    1000101100101111    1000101100110000    1000101100110001    1000101100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35630 - 35634

  --1000101100110011    1000101100110100    1000101100110101    1000101100110110    1000101100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35635 - 35639

  --1000101100111000    1000101100111001    1000101100111010    1000101100111011    1000101100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35640 - 35644

  --1000101100111101    1000101100111110    1000101100111111    1000101101000000    1000101101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35645 - 35649

  --1000101101000010    1000101101000011    1000101101000100    1000101101000101    1000101101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35650 - 35654

  --1000101101000111    1000101101001000    1000101101001001    1000101101001010    1000101101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35655 - 35659

  --1000101101001100    1000101101001101    1000101101001110    1000101101001111    1000101101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35660 - 35664

  --1000101101010001    1000101101010010    1000101101010011    1000101101010100    1000101101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35665 - 35669

  --1000101101010110    1000101101010111    1000101101011000    1000101101011001    1000101101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35670 - 35674

  --1000101101011011    1000101101011100    1000101101011101    1000101101011110    1000101101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35675 - 35679

  --1000101101100000    1000101101100001    1000101101100010    1000101101100011    1000101101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35680 - 35684

  --1000101101100101    1000101101100110    1000101101100111    1000101101101000    1000101101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35685 - 35689

  --1000101101101010    1000101101101011    1000101101101100    1000101101101101    1000101101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35690 - 35694

  --1000101101101111    1000101101110000    1000101101110001    1000101101110010    1000101101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35695 - 35699

  --1000101101110100    1000101101110101    1000101101110110    1000101101110111    1000101101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35700 - 35704

  --1000101101111001    1000101101111010    1000101101111011    1000101101111100    1000101101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35705 - 35709

  --1000101101111110    1000101101111111    1000101110000000    1000101110000001    1000101110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35710 - 35714

  --1000101110000011    1000101110000100    1000101110000101    1000101110000110    1000101110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35715 - 35719

  --1000101110001000    1000101110001001    1000101110001010    1000101110001011    1000101110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35720 - 35724

  --1000101110001101    1000101110001110    1000101110001111    1000101110010000    1000101110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35725 - 35729

  --1000101110010010    1000101110010011    1000101110010100    1000101110010101    1000101110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35730 - 35734

  --1000101110010111    1000101110011000    1000101110011001    1000101110011010    1000101110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35735 - 35739

  --1000101110011100    1000101110011101    1000101110011110    1000101110011111    1000101110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35740 - 35744

  --1000101110100001    1000101110100010    1000101110100011    1000101110100100    1000101110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35745 - 35749

  --1000101110100110    1000101110100111    1000101110101000    1000101110101001    1000101110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35750 - 35754

  --1000101110101011    1000101110101100    1000101110101101    1000101110101110    1000101110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35755 - 35759

  --1000101110110000    1000101110110001    1000101110110010    1000101110110011    1000101110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35760 - 35764

  --1000101110110101    1000101110110110    1000101110110111    1000101110111000    1000101110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35765 - 35769

  --1000101110111010    1000101110111011    1000101110111100    1000101110111101    1000101110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35770 - 35774

  --1000101110111111    1000101111000000    1000101111000001    1000101111000010    1000101111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35775 - 35779

  --1000101111000100    1000101111000101    1000101111000110    1000101111000111    1000101111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35780 - 35784

  --1000101111001001    1000101111001010    1000101111001011    1000101111001100    1000101111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35785 - 35789

  --1000101111001110    1000101111001111    1000101111010000    1000101111010001    1000101111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35790 - 35794

  --1000101111010011    1000101111010100    1000101111010101    1000101111010110    1000101111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35795 - 35799

  --1000101111011000    1000101111011001    1000101111011010    1000101111011011    1000101111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35800 - 35804

  --1000101111011101    1000101111011110    1000101111011111    1000101111100000    1000101111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35805 - 35809

  --1000101111100010    1000101111100011    1000101111100100    1000101111100101    1000101111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35810 - 35814

  --1000101111100111    1000101111101000    1000101111101001    1000101111101010    1000101111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35815 - 35819

  --1000101111101100    1000101111101101    1000101111101110    1000101111101111    1000101111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35820 - 35824

  --1000101111110001    1000101111110010    1000101111110011    1000101111110100    1000101111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35825 - 35829

  --1000101111110110    1000101111110111    1000101111111000    1000101111111001    1000101111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35830 - 35834

  --1000101111111011    1000101111111100    1000101111111101    1000101111111110    1000101111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35835 - 35839

  --1000110000000000    1000110000000001    1000110000000010    1000110000000011    1000110000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35840 - 35844

  --1000110000000101    1000110000000110    1000110000000111    1000110000001000    1000110000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35845 - 35849

  --1000110000001010    1000110000001011    1000110000001100    1000110000001101    1000110000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35850 - 35854

  --1000110000001111    1000110000010000    1000110000010001    1000110000010010    1000110000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35855 - 35859

  --1000110000010100    1000110000010101    1000110000010110    1000110000010111    1000110000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35860 - 35864

  --1000110000011001    1000110000011010    1000110000011011    1000110000011100    1000110000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35865 - 35869

  --1000110000011110    1000110000011111    1000110000100000    1000110000100001    1000110000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35870 - 35874

  --1000110000100011    1000110000100100    1000110000100101    1000110000100110    1000110000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35875 - 35879

  --1000110000101000    1000110000101001    1000110000101010    1000110000101011    1000110000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35880 - 35884

  --1000110000101101    1000110000101110    1000110000101111    1000110000110000    1000110000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35885 - 35889

  --1000110000110010    1000110000110011    1000110000110100    1000110000110101    1000110000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35890 - 35894

  --1000110000110111    1000110000111000    1000110000111001    1000110000111010    1000110000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35895 - 35899

  --1000110000111100    1000110000111101    1000110000111110    1000110000111111    1000110001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35900 - 35904

  --1000110001000001    1000110001000010    1000110001000011    1000110001000100    1000110001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35905 - 35909

  --1000110001000110    1000110001000111    1000110001001000    1000110001001001    1000110001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35910 - 35914

  --1000110001001011    1000110001001100    1000110001001101    1000110001001110    1000110001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35915 - 35919

  --1000110001010000    1000110001010001    1000110001010010    1000110001010011    1000110001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35920 - 35924

  --1000110001010101    1000110001010110    1000110001010111    1000110001011000    1000110001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35925 - 35929

  --1000110001011010    1000110001011011    1000110001011100    1000110001011101    1000110001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35930 - 35934

  --1000110001011111    1000110001100000    1000110001100001    1000110001100010    1000110001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35935 - 35939

  --1000110001100100    1000110001100101    1000110001100110    1000110001100111    1000110001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35940 - 35944

  --1000110001101001    1000110001101010    1000110001101011    1000110001101100    1000110001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35945 - 35949

  --1000110001101110    1000110001101111    1000110001110000    1000110001110001    1000110001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35950 - 35954

  --1000110001110011    1000110001110100    1000110001110101    1000110001110110    1000110001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35955 - 35959

  --1000110001111000    1000110001111001    1000110001111010    1000110001111011    1000110001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35960 - 35964

  --1000110001111101    1000110001111110    1000110001111111    1000110010000000    1000110010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35965 - 35969

  --1000110010000010    1000110010000011    1000110010000100    1000110010000101    1000110010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35970 - 35974

  --1000110010000111    1000110010001000    1000110010001001    1000110010001010    1000110010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35975 - 35979

  --1000110010001100    1000110010001101    1000110010001110    1000110010001111    1000110010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35980 - 35984

  --1000110010010001    1000110010010010    1000110010010011    1000110010010100    1000110010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35985 - 35989

  --1000110010010110    1000110010010111    1000110010011000    1000110010011001    1000110010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35990 - 35994

  --1000110010011011    1000110010011100    1000110010011101    1000110010011110    1000110010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 35995 - 35999

  --1000110010100000    1000110010100001    1000110010100010    1000110010100011    1000110010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36000 - 36004

  --1000110010100101    1000110010100110    1000110010100111    1000110010101000    1000110010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36005 - 36009

  --1000110010101010    1000110010101011    1000110010101100    1000110010101101    1000110010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36010 - 36014

  --1000110010101111    1000110010110000    1000110010110001    1000110010110010    1000110010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36015 - 36019

  --1000110010110100    1000110010110101    1000110010110110    1000110010110111    1000110010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36020 - 36024

  --1000110010111001    1000110010111010    1000110010111011    1000110010111100    1000110010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36025 - 36029

  --1000110010111110    1000110010111111    1000110011000000    1000110011000001    1000110011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36030 - 36034

  --1000110011000011    1000110011000100    1000110011000101    1000110011000110    1000110011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36035 - 36039

  --1000110011001000    1000110011001001    1000110011001010    1000110011001011    1000110011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36040 - 36044

  --1000110011001101    1000110011001110    1000110011001111    1000110011010000    1000110011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36045 - 36049

  --1000110011010010    1000110011010011    1000110011010100    1000110011010101    1000110011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36050 - 36054

  --1000110011010111    1000110011011000    1000110011011001    1000110011011010    1000110011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36055 - 36059

  --1000110011011100    1000110011011101    1000110011011110    1000110011011111    1000110011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36060 - 36064

  --1000110011100001    1000110011100010    1000110011100011    1000110011100100    1000110011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36065 - 36069

  --1000110011100110    1000110011100111    1000110011101000    1000110011101001    1000110011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36070 - 36074

  --1000110011101011    1000110011101100    1000110011101101    1000110011101110    1000110011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36075 - 36079

  --1000110011110000    1000110011110001    1000110011110010    1000110011110011    1000110011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36080 - 36084

  --1000110011110101    1000110011110110    1000110011110111    1000110011111000    1000110011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36085 - 36089

  --1000110011111010    1000110011111011    1000110011111100    1000110011111101    1000110011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36090 - 36094

  --1000110011111111    1000110100000000    1000110100000001    1000110100000010    1000110100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36095 - 36099

  --1000110100000100    1000110100000101    1000110100000110    1000110100000111    1000110100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36100 - 36104

  --1000110100001001    1000110100001010    1000110100001011    1000110100001100    1000110100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36105 - 36109

  --1000110100001110    1000110100001111    1000110100010000    1000110100010001    1000110100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36110 - 36114

  --1000110100010011    1000110100010100    1000110100010101    1000110100010110    1000110100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36115 - 36119

  --1000110100011000    1000110100011001    1000110100011010    1000110100011011    1000110100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36120 - 36124

  --1000110100011101    1000110100011110    1000110100011111    1000110100100000    1000110100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36125 - 36129

  --1000110100100010    1000110100100011    1000110100100100    1000110100100101    1000110100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36130 - 36134

  --1000110100100111    1000110100101000    1000110100101001    1000110100101010    1000110100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36135 - 36139

  --1000110100101100    1000110100101101    1000110100101110    1000110100101111    1000110100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36140 - 36144

  --1000110100110001    1000110100110010    1000110100110011    1000110100110100    1000110100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36145 - 36149

  --1000110100110110    1000110100110111    1000110100111000    1000110100111001    1000110100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36150 - 36154

  --1000110100111011    1000110100111100    1000110100111101    1000110100111110    1000110100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36155 - 36159

  --1000110101000000    1000110101000001    1000110101000010    1000110101000011    1000110101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36160 - 36164

  --1000110101000101    1000110101000110    1000110101000111    1000110101001000    1000110101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36165 - 36169

  --1000110101001010    1000110101001011    1000110101001100    1000110101001101    1000110101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36170 - 36174

  --1000110101001111    1000110101010000    1000110101010001    1000110101010010    1000110101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36175 - 36179

  --1000110101010100    1000110101010101    1000110101010110    1000110101010111    1000110101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36180 - 36184

  --1000110101011001    1000110101011010    1000110101011011    1000110101011100    1000110101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36185 - 36189

  --1000110101011110    1000110101011111    1000110101100000    1000110101100001    1000110101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36190 - 36194

  --1000110101100011    1000110101100100    1000110101100101    1000110101100110    1000110101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36195 - 36199

  --1000110101101000    1000110101101001    1000110101101010    1000110101101011    1000110101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36200 - 36204

  --1000110101101101    1000110101101110    1000110101101111    1000110101110000    1000110101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36205 - 36209

  --1000110101110010    1000110101110011    1000110101110100    1000110101110101    1000110101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36210 - 36214

  --1000110101110111    1000110101111000    1000110101111001    1000110101111010    1000110101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36215 - 36219

  --1000110101111100    1000110101111101    1000110101111110    1000110101111111    1000110110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36220 - 36224

  --1000110110000001    1000110110000010    1000110110000011    1000110110000100    1000110110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36225 - 36229

  --1000110110000110    1000110110000111    1000110110001000    1000110110001001    1000110110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36230 - 36234

  --1000110110001011    1000110110001100    1000110110001101    1000110110001110    1000110110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36235 - 36239

  --1000110110010000    1000110110010001    1000110110010010    1000110110010011    1000110110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36240 - 36244

  --1000110110010101    1000110110010110    1000110110010111    1000110110011000    1000110110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36245 - 36249

  --1000110110011010    1000110110011011    1000110110011100    1000110110011101    1000110110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36250 - 36254

  --1000110110011111    1000110110100000    1000110110100001    1000110110100010    1000110110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36255 - 36259

  --1000110110100100    1000110110100101    1000110110100110    1000110110100111    1000110110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36260 - 36264

  --1000110110101001    1000110110101010    1000110110101011    1000110110101100    1000110110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36265 - 36269

  --1000110110101110    1000110110101111    1000110110110000    1000110110110001    1000110110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36270 - 36274

  --1000110110110011    1000110110110100    1000110110110101    1000110110110110    1000110110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36275 - 36279

  --1000110110111000    1000110110111001    1000110110111010    1000110110111011    1000110110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36280 - 36284

  --1000110110111101    1000110110111110    1000110110111111    1000110111000000    1000110111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36285 - 36289

  --1000110111000010    1000110111000011    1000110111000100    1000110111000101    1000110111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36290 - 36294

  --1000110111000111    1000110111001000    1000110111001001    1000110111001010    1000110111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36295 - 36299

  --1000110111001100    1000110111001101    1000110111001110    1000110111001111    1000110111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36300 - 36304

  --1000110111010001    1000110111010010    1000110111010011    1000110111010100    1000110111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36305 - 36309

  --1000110111010110    1000110111010111    1000110111011000    1000110111011001    1000110111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36310 - 36314

  --1000110111011011    1000110111011100    1000110111011101    1000110111011110    1000110111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36315 - 36319

  --1000110111100000    1000110111100001    1000110111100010    1000110111100011    1000110111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36320 - 36324

  --1000110111100101    1000110111100110    1000110111100111    1000110111101000    1000110111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36325 - 36329

  --1000110111101010    1000110111101011    1000110111101100    1000110111101101    1000110111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36330 - 36334

  --1000110111101111    1000110111110000    1000110111110001    1000110111110010    1000110111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36335 - 36339

  --1000110111110100    1000110111110101    1000110111110110    1000110111110111    1000110111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36340 - 36344

  --1000110111111001    1000110111111010    1000110111111011    1000110111111100    1000110111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36345 - 36349

  --1000110111111110    1000110111111111    1000111000000000    1000111000000001    1000111000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36350 - 36354

  --1000111000000011    1000111000000100    1000111000000101    1000111000000110    1000111000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36355 - 36359

  --1000111000001000    1000111000001001    1000111000001010    1000111000001011    1000111000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36360 - 36364

  --1000111000001101    1000111000001110    1000111000001111    1000111000010000    1000111000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36365 - 36369

  --1000111000010010    1000111000010011    1000111000010100    1000111000010101    1000111000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36370 - 36374

  --1000111000010111    1000111000011000    1000111000011001    1000111000011010    1000111000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36375 - 36379

  --1000111000011100    1000111000011101    1000111000011110    1000111000011111    1000111000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36380 - 36384

  --1000111000100001    1000111000100010    1000111000100011    1000111000100100    1000111000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36385 - 36389

  --1000111000100110    1000111000100111    1000111000101000    1000111000101001    1000111000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36390 - 36394

  --1000111000101011    1000111000101100    1000111000101101    1000111000101110    1000111000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36395 - 36399

  --1000111000110000    1000111000110001    1000111000110010    1000111000110011    1000111000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36400 - 36404

  --1000111000110101    1000111000110110    1000111000110111    1000111000111000    1000111000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36405 - 36409

  --1000111000111010    1000111000111011    1000111000111100    1000111000111101    1000111000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36410 - 36414

  --1000111000111111    1000111001000000    1000111001000001    1000111001000010    1000111001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36415 - 36419

  --1000111001000100    1000111001000101    1000111001000110    1000111001000111    1000111001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36420 - 36424

  --1000111001001001    1000111001001010    1000111001001011    1000111001001100    1000111001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36425 - 36429

  --1000111001001110    1000111001001111    1000111001010000    1000111001010001    1000111001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36430 - 36434

  --1000111001010011    1000111001010100    1000111001010101    1000111001010110    1000111001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36435 - 36439

  --1000111001011000    1000111001011001    1000111001011010    1000111001011011    1000111001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36440 - 36444

  --1000111001011101    1000111001011110    1000111001011111    1000111001100000    1000111001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36445 - 36449

  --1000111001100010    1000111001100011    1000111001100100    1000111001100101    1000111001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36450 - 36454

  --1000111001100111    1000111001101000    1000111001101001    1000111001101010    1000111001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36455 - 36459

  --1000111001101100    1000111001101101    1000111001101110    1000111001101111    1000111001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36460 - 36464

  --1000111001110001    1000111001110010    1000111001110011    1000111001110100    1000111001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36465 - 36469

  --1000111001110110    1000111001110111    1000111001111000    1000111001111001    1000111001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36470 - 36474

  --1000111001111011    1000111001111100    1000111001111101    1000111001111110    1000111001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36475 - 36479

  --1000111010000000    1000111010000001    1000111010000010    1000111010000011    1000111010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36480 - 36484

  --1000111010000101    1000111010000110    1000111010000111    1000111010001000    1000111010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36485 - 36489

  --1000111010001010    1000111010001011    1000111010001100    1000111010001101    1000111010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36490 - 36494

  --1000111010001111    1000111010010000    1000111010010001    1000111010010010    1000111010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36495 - 36499

  --1000111010010100    1000111010010101    1000111010010110    1000111010010111    1000111010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36500 - 36504

  --1000111010011001    1000111010011010    1000111010011011    1000111010011100    1000111010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36505 - 36509

  --1000111010011110    1000111010011111    1000111010100000    1000111010100001    1000111010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36510 - 36514

  --1000111010100011    1000111010100100    1000111010100101    1000111010100110    1000111010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36515 - 36519

  --1000111010101000    1000111010101001    1000111010101010    1000111010101011    1000111010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36520 - 36524

  --1000111010101101    1000111010101110    1000111010101111    1000111010110000    1000111010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36525 - 36529

  --1000111010110010    1000111010110011    1000111010110100    1000111010110101    1000111010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36530 - 36534

  --1000111010110111    1000111010111000    1000111010111001    1000111010111010    1000111010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36535 - 36539

  --1000111010111100    1000111010111101    1000111010111110    1000111010111111    1000111011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36540 - 36544

  --1000111011000001    1000111011000010    1000111011000011    1000111011000100    1000111011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36545 - 36549

  --1000111011000110    1000111011000111    1000111011001000    1000111011001001    1000111011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36550 - 36554

  --1000111011001011    1000111011001100    1000111011001101    1000111011001110    1000111011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36555 - 36559

  --1000111011010000    1000111011010001    1000111011010010    1000111011010011    1000111011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36560 - 36564

  --1000111011010101    1000111011010110    1000111011010111    1000111011011000    1000111011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36565 - 36569

  --1000111011011010    1000111011011011    1000111011011100    1000111011011101    1000111011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36570 - 36574

  --1000111011011111    1000111011100000    1000111011100001    1000111011100010    1000111011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36575 - 36579

  --1000111011100100    1000111011100101    1000111011100110    1000111011100111    1000111011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36580 - 36584

  --1000111011101001    1000111011101010    1000111011101011    1000111011101100    1000111011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36585 - 36589

  --1000111011101110    1000111011101111    1000111011110000    1000111011110001    1000111011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36590 - 36594

  --1000111011110011    1000111011110100    1000111011110101    1000111011110110    1000111011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36595 - 36599

  --1000111011111000    1000111011111001    1000111011111010    1000111011111011    1000111011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36600 - 36604

  --1000111011111101    1000111011111110    1000111011111111    1000111100000000    1000111100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36605 - 36609

  --1000111100000010    1000111100000011    1000111100000100    1000111100000101    1000111100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36610 - 36614

  --1000111100000111    1000111100001000    1000111100001001    1000111100001010    1000111100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36615 - 36619

  --1000111100001100    1000111100001101    1000111100001110    1000111100001111    1000111100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36620 - 36624

  --1000111100010001    1000111100010010    1000111100010011    1000111100010100    1000111100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36625 - 36629

  --1000111100010110    1000111100010111    1000111100011000    1000111100011001    1000111100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36630 - 36634

  --1000111100011011    1000111100011100    1000111100011101    1000111100011110    1000111100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36635 - 36639

  --1000111100100000    1000111100100001    1000111100100010    1000111100100011    1000111100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36640 - 36644

  --1000111100100101    1000111100100110    1000111100100111    1000111100101000    1000111100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36645 - 36649

  --1000111100101010    1000111100101011    1000111100101100    1000111100101101    1000111100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36650 - 36654

  --1000111100101111    1000111100110000    1000111100110001    1000111100110010    1000111100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36655 - 36659

  --1000111100110100    1000111100110101    1000111100110110    1000111100110111    1000111100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36660 - 36664

  --1000111100111001    1000111100111010    1000111100111011    1000111100111100    1000111100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36665 - 36669

  --1000111100111110    1000111100111111    1000111101000000    1000111101000001    1000111101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36670 - 36674

  --1000111101000011    1000111101000100    1000111101000101    1000111101000110    1000111101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36675 - 36679

  --1000111101001000    1000111101001001    1000111101001010    1000111101001011    1000111101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36680 - 36684

  --1000111101001101    1000111101001110    1000111101001111    1000111101010000    1000111101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36685 - 36689

  --1000111101010010    1000111101010011    1000111101010100    1000111101010101    1000111101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36690 - 36694

  --1000111101010111    1000111101011000    1000111101011001    1000111101011010    1000111101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36695 - 36699

  --1000111101011100    1000111101011101    1000111101011110    1000111101011111    1000111101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36700 - 36704

  --1000111101100001    1000111101100010    1000111101100011    1000111101100100    1000111101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36705 - 36709

  --1000111101100110    1000111101100111    1000111101101000    1000111101101001    1000111101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36710 - 36714

  --1000111101101011    1000111101101100    1000111101101101    1000111101101110    1000111101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36715 - 36719

  --1000111101110000    1000111101110001    1000111101110010    1000111101110011    1000111101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36720 - 36724

  --1000111101110101    1000111101110110    1000111101110111    1000111101111000    1000111101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36725 - 36729

  --1000111101111010    1000111101111011    1000111101111100    1000111101111101    1000111101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36730 - 36734

  --1000111101111111    1000111110000000    1000111110000001    1000111110000010    1000111110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36735 - 36739

  --1000111110000100    1000111110000101    1000111110000110    1000111110000111    1000111110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36740 - 36744

  --1000111110001001    1000111110001010    1000111110001011    1000111110001100    1000111110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36745 - 36749

  --1000111110001110    1000111110001111    1000111110010000    1000111110010001    1000111110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36750 - 36754

  --1000111110010011    1000111110010100    1000111110010101    1000111110010110    1000111110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36755 - 36759

  --1000111110011000    1000111110011001    1000111110011010    1000111110011011    1000111110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36760 - 36764

  --1000111110011101    1000111110011110    1000111110011111    1000111110100000    1000111110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36765 - 36769

  --1000111110100010    1000111110100011    1000111110100100    1000111110100101    1000111110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36770 - 36774

  --1000111110100111    1000111110101000    1000111110101001    1000111110101010    1000111110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36775 - 36779

  --1000111110101100    1000111110101101    1000111110101110    1000111110101111    1000111110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36780 - 36784

  --1000111110110001    1000111110110010    1000111110110011    1000111110110100    1000111110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36785 - 36789

  --1000111110110110    1000111110110111    1000111110111000    1000111110111001    1000111110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36790 - 36794

  --1000111110111011    1000111110111100    1000111110111101    1000111110111110    1000111110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36795 - 36799

  --1000111111000000    1000111111000001    1000111111000010    1000111111000011    1000111111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36800 - 36804

  --1000111111000101    1000111111000110    1000111111000111    1000111111001000    1000111111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36805 - 36809

  --1000111111001010    1000111111001011    1000111111001100    1000111111001101    1000111111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36810 - 36814

  --1000111111001111    1000111111010000    1000111111010001    1000111111010010    1000111111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36815 - 36819

  --1000111111010100    1000111111010101    1000111111010110    1000111111010111    1000111111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36820 - 36824

  --1000111111011001    1000111111011010    1000111111011011    1000111111011100    1000111111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36825 - 36829

  --1000111111011110    1000111111011111    1000111111100000    1000111111100001    1000111111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36830 - 36834

  --1000111111100011    1000111111100100    1000111111100101    1000111111100110    1000111111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36835 - 36839

  --1000111111101000    1000111111101001    1000111111101010    1000111111101011    1000111111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36840 - 36844

  --1000111111101101    1000111111101110    1000111111101111    1000111111110000    1000111111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36845 - 36849

  --1000111111110010    1000111111110011    1000111111110100    1000111111110101    1000111111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36850 - 36854

  --1000111111110111    1000111111111000    1000111111111001    1000111111111010    1000111111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36855 - 36859

  --1000111111111100    1000111111111101    1000111111111110    1000111111111111    1001000000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36860 - 36864

  --1001000000000001    1001000000000010    1001000000000011    1001000000000100    1001000000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36865 - 36869

  --1001000000000110    1001000000000111    1001000000001000    1001000000001001    1001000000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36870 - 36874

  --1001000000001011    1001000000001100    1001000000001101    1001000000001110    1001000000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36875 - 36879

  --1001000000010000    1001000000010001    1001000000010010    1001000000010011    1001000000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36880 - 36884

  --1001000000010101    1001000000010110    1001000000010111    1001000000011000    1001000000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36885 - 36889

  --1001000000011010    1001000000011011    1001000000011100    1001000000011101    1001000000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36890 - 36894

  --1001000000011111    1001000000100000    1001000000100001    1001000000100010    1001000000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36895 - 36899

  --1001000000100100    1001000000100101    1001000000100110    1001000000100111    1001000000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36900 - 36904

  --1001000000101001    1001000000101010    1001000000101011    1001000000101100    1001000000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36905 - 36909

  --1001000000101110    1001000000101111    1001000000110000    1001000000110001    1001000000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36910 - 36914

  --1001000000110011    1001000000110100    1001000000110101    1001000000110110    1001000000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36915 - 36919

  --1001000000111000    1001000000111001    1001000000111010    1001000000111011    1001000000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36920 - 36924

  --1001000000111101    1001000000111110    1001000000111111    1001000001000000    1001000001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36925 - 36929

  --1001000001000010    1001000001000011    1001000001000100    1001000001000101    1001000001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36930 - 36934

  --1001000001000111    1001000001001000    1001000001001001    1001000001001010    1001000001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36935 - 36939

  --1001000001001100    1001000001001101    1001000001001110    1001000001001111    1001000001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36940 - 36944

  --1001000001010001    1001000001010010    1001000001010011    1001000001010100    1001000001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36945 - 36949

  --1001000001010110    1001000001010111    1001000001011000    1001000001011001    1001000001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36950 - 36954

  --1001000001011011    1001000001011100    1001000001011101    1001000001011110    1001000001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36955 - 36959

  --1001000001100000    1001000001100001    1001000001100010    1001000001100011    1001000001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36960 - 36964

  --1001000001100101    1001000001100110    1001000001100111    1001000001101000    1001000001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36965 - 36969

  --1001000001101010    1001000001101011    1001000001101100    1001000001101101    1001000001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36970 - 36974

  --1001000001101111    1001000001110000    1001000001110001    1001000001110010    1001000001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36975 - 36979

  --1001000001110100    1001000001110101    1001000001110110    1001000001110111    1001000001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36980 - 36984

  --1001000001111001    1001000001111010    1001000001111011    1001000001111100    1001000001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36985 - 36989

  --1001000001111110    1001000001111111    1001000010000000    1001000010000001    1001000010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36990 - 36994

  --1001000010000011    1001000010000100    1001000010000101    1001000010000110    1001000010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 36995 - 36999

  --1001000010001000    1001000010001001    1001000010001010    1001000010001011    1001000010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37000 - 37004

  --1001000010001101    1001000010001110    1001000010001111    1001000010010000    1001000010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37005 - 37009

  --1001000010010010    1001000010010011    1001000010010100    1001000010010101    1001000010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37010 - 37014

  --1001000010010111    1001000010011000    1001000010011001    1001000010011010    1001000010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37015 - 37019

  --1001000010011100    1001000010011101    1001000010011110    1001000010011111    1001000010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37020 - 37024

  --1001000010100001    1001000010100010    1001000010100011    1001000010100100    1001000010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37025 - 37029

  --1001000010100110    1001000010100111    1001000010101000    1001000010101001    1001000010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37030 - 37034

  --1001000010101011    1001000010101100    1001000010101101    1001000010101110    1001000010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37035 - 37039

  --1001000010110000    1001000010110001    1001000010110010    1001000010110011    1001000010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37040 - 37044

  --1001000010110101    1001000010110110    1001000010110111    1001000010111000    1001000010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37045 - 37049

  --1001000010111010    1001000010111011    1001000010111100    1001000010111101    1001000010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37050 - 37054

  --1001000010111111    1001000011000000    1001000011000001    1001000011000010    1001000011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37055 - 37059

  --1001000011000100    1001000011000101    1001000011000110    1001000011000111    1001000011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37060 - 37064

  --1001000011001001    1001000011001010    1001000011001011    1001000011001100    1001000011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37065 - 37069

  --1001000011001110    1001000011001111    1001000011010000    1001000011010001    1001000011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37070 - 37074

  --1001000011010011    1001000011010100    1001000011010101    1001000011010110    1001000011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37075 - 37079

  --1001000011011000    1001000011011001    1001000011011010    1001000011011011    1001000011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37080 - 37084

  --1001000011011101    1001000011011110    1001000011011111    1001000011100000    1001000011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37085 - 37089

  --1001000011100010    1001000011100011    1001000011100100    1001000011100101    1001000011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37090 - 37094

  --1001000011100111    1001000011101000    1001000011101001    1001000011101010    1001000011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37095 - 37099

  --1001000011101100    1001000011101101    1001000011101110    1001000011101111    1001000011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37100 - 37104

  --1001000011110001    1001000011110010    1001000011110011    1001000011110100    1001000011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37105 - 37109

  --1001000011110110    1001000011110111    1001000011111000    1001000011111001    1001000011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37110 - 37114

  --1001000011111011    1001000011111100    1001000011111101    1001000011111110    1001000011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37115 - 37119

  --1001000100000000    1001000100000001    1001000100000010    1001000100000011    1001000100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37120 - 37124

  --1001000100000101    1001000100000110    1001000100000111    1001000100001000    1001000100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37125 - 37129

  --1001000100001010    1001000100001011    1001000100001100    1001000100001101    1001000100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37130 - 37134

  --1001000100001111    1001000100010000    1001000100010001    1001000100010010    1001000100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37135 - 37139

  --1001000100010100    1001000100010101    1001000100010110    1001000100010111    1001000100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37140 - 37144

  --1001000100011001    1001000100011010    1001000100011011    1001000100011100    1001000100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37145 - 37149

  --1001000100011110    1001000100011111    1001000100100000    1001000100100001    1001000100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37150 - 37154

  --1001000100100011    1001000100100100    1001000100100101    1001000100100110    1001000100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37155 - 37159

  --1001000100101000    1001000100101001    1001000100101010    1001000100101011    1001000100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37160 - 37164

  --1001000100101101    1001000100101110    1001000100101111    1001000100110000    1001000100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37165 - 37169

  --1001000100110010    1001000100110011    1001000100110100    1001000100110101    1001000100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37170 - 37174

  --1001000100110111    1001000100111000    1001000100111001    1001000100111010    1001000100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37175 - 37179

  --1001000100111100    1001000100111101    1001000100111110    1001000100111111    1001000101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37180 - 37184

  --1001000101000001    1001000101000010    1001000101000011    1001000101000100    1001000101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37185 - 37189

  --1001000101000110    1001000101000111    1001000101001000    1001000101001001    1001000101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37190 - 37194

  --1001000101001011    1001000101001100    1001000101001101    1001000101001110    1001000101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37195 - 37199

  --1001000101010000    1001000101010001    1001000101010010    1001000101010011    1001000101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37200 - 37204

  --1001000101010101    1001000101010110    1001000101010111    1001000101011000    1001000101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37205 - 37209

  --1001000101011010    1001000101011011    1001000101011100    1001000101011101    1001000101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37210 - 37214

  --1001000101011111    1001000101100000    1001000101100001    1001000101100010    1001000101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37215 - 37219

  --1001000101100100    1001000101100101    1001000101100110    1001000101100111    1001000101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37220 - 37224

  --1001000101101001    1001000101101010    1001000101101011    1001000101101100    1001000101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37225 - 37229

  --1001000101101110    1001000101101111    1001000101110000    1001000101110001    1001000101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37230 - 37234

  --1001000101110011    1001000101110100    1001000101110101    1001000101110110    1001000101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37235 - 37239

  --1001000101111000    1001000101111001    1001000101111010    1001000101111011    1001000101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37240 - 37244

  --1001000101111101    1001000101111110    1001000101111111    1001000110000000    1001000110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37245 - 37249

  --1001000110000010    1001000110000011    1001000110000100    1001000110000101    1001000110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37250 - 37254

  --1001000110000111    1001000110001000    1001000110001001    1001000110001010    1001000110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37255 - 37259

  --1001000110001100    1001000110001101    1001000110001110    1001000110001111    1001000110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37260 - 37264

  --1001000110010001    1001000110010010    1001000110010011    1001000110010100    1001000110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37265 - 37269

  --1001000110010110    1001000110010111    1001000110011000    1001000110011001    1001000110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37270 - 37274

  --1001000110011011    1001000110011100    1001000110011101    1001000110011110    1001000110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37275 - 37279

  --1001000110100000    1001000110100001    1001000110100010    1001000110100011    1001000110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37280 - 37284

  --1001000110100101    1001000110100110    1001000110100111    1001000110101000    1001000110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37285 - 37289

  --1001000110101010    1001000110101011    1001000110101100    1001000110101101    1001000110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37290 - 37294

  --1001000110101111    1001000110110000    1001000110110001    1001000110110010    1001000110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37295 - 37299

  --1001000110110100    1001000110110101    1001000110110110    1001000110110111    1001000110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37300 - 37304

  --1001000110111001    1001000110111010    1001000110111011    1001000110111100    1001000110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37305 - 37309

  --1001000110111110    1001000110111111    1001000111000000    1001000111000001    1001000111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37310 - 37314

  --1001000111000011    1001000111000100    1001000111000101    1001000111000110    1001000111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37315 - 37319

  --1001000111001000    1001000111001001    1001000111001010    1001000111001011    1001000111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37320 - 37324

  --1001000111001101    1001000111001110    1001000111001111    1001000111010000    1001000111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37325 - 37329

  --1001000111010010    1001000111010011    1001000111010100    1001000111010101    1001000111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37330 - 37334

  --1001000111010111    1001000111011000    1001000111011001    1001000111011010    1001000111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37335 - 37339

  --1001000111011100    1001000111011101    1001000111011110    1001000111011111    1001000111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37340 - 37344

  --1001000111100001    1001000111100010    1001000111100011    1001000111100100    1001000111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37345 - 37349

  --1001000111100110    1001000111100111    1001000111101000    1001000111101001    1001000111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37350 - 37354

  --1001000111101011    1001000111101100    1001000111101101    1001000111101110    1001000111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37355 - 37359

  --1001000111110000    1001000111110001    1001000111110010    1001000111110011    1001000111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37360 - 37364

  --1001000111110101    1001000111110110    1001000111110111    1001000111111000    1001000111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37365 - 37369

  --1001000111111010    1001000111111011    1001000111111100    1001000111111101    1001000111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37370 - 37374

  --1001000111111111    1001001000000000    1001001000000001    1001001000000010    1001001000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37375 - 37379

  --1001001000000100    1001001000000101    1001001000000110    1001001000000111    1001001000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37380 - 37384

  --1001001000001001    1001001000001010    1001001000001011    1001001000001100    1001001000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37385 - 37389

  --1001001000001110    1001001000001111    1001001000010000    1001001000010001    1001001000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37390 - 37394

  --1001001000010011    1001001000010100    1001001000010101    1001001000010110    1001001000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37395 - 37399

  --1001001000011000    1001001000011001    1001001000011010    1001001000011011    1001001000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37400 - 37404

  --1001001000011101    1001001000011110    1001001000011111    1001001000100000    1001001000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37405 - 37409

  --1001001000100010    1001001000100011    1001001000100100    1001001000100101    1001001000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37410 - 37414

  --1001001000100111    1001001000101000    1001001000101001    1001001000101010    1001001000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37415 - 37419

  --1001001000101100    1001001000101101    1001001000101110    1001001000101111    1001001000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37420 - 37424

  --1001001000110001    1001001000110010    1001001000110011    1001001000110100    1001001000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37425 - 37429

  --1001001000110110    1001001000110111    1001001000111000    1001001000111001    1001001000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37430 - 37434

  --1001001000111011    1001001000111100    1001001000111101    1001001000111110    1001001000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37435 - 37439

  --1001001001000000    1001001001000001    1001001001000010    1001001001000011    1001001001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37440 - 37444

  --1001001001000101    1001001001000110    1001001001000111    1001001001001000    1001001001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37445 - 37449

  --1001001001001010    1001001001001011    1001001001001100    1001001001001101    1001001001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37450 - 37454

  --1001001001001111    1001001001010000    1001001001010001    1001001001010010    1001001001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37455 - 37459

  --1001001001010100    1001001001010101    1001001001010110    1001001001010111    1001001001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37460 - 37464

  --1001001001011001    1001001001011010    1001001001011011    1001001001011100    1001001001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37465 - 37469

  --1001001001011110    1001001001011111    1001001001100000    1001001001100001    1001001001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37470 - 37474

  --1001001001100011    1001001001100100    1001001001100101    1001001001100110    1001001001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37475 - 37479

  --1001001001101000    1001001001101001    1001001001101010    1001001001101011    1001001001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37480 - 37484

  --1001001001101101    1001001001101110    1001001001101111    1001001001110000    1001001001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37485 - 37489

  --1001001001110010    1001001001110011    1001001001110100    1001001001110101    1001001001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37490 - 37494

  --1001001001110111    1001001001111000    1001001001111001    1001001001111010    1001001001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37495 - 37499

  --1001001001111100    1001001001111101    1001001001111110    1001001001111111    1001001010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37500 - 37504

  --1001001010000001    1001001010000010    1001001010000011    1001001010000100    1001001010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37505 - 37509

  --1001001010000110    1001001010000111    1001001010001000    1001001010001001    1001001010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37510 - 37514

  --1001001010001011    1001001010001100    1001001010001101    1001001010001110    1001001010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37515 - 37519

  --1001001010010000    1001001010010001    1001001010010010    1001001010010011    1001001010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37520 - 37524

  --1001001010010101    1001001010010110    1001001010010111    1001001010011000    1001001010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37525 - 37529

  --1001001010011010    1001001010011011    1001001010011100    1001001010011101    1001001010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37530 - 37534

  --1001001010011111    1001001010100000    1001001010100001    1001001010100010    1001001010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37535 - 37539

  --1001001010100100    1001001010100101    1001001010100110    1001001010100111    1001001010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37540 - 37544

  --1001001010101001    1001001010101010    1001001010101011    1001001010101100    1001001010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37545 - 37549

  --1001001010101110    1001001010101111    1001001010110000    1001001010110001    1001001010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37550 - 37554

  --1001001010110011    1001001010110100    1001001010110101    1001001010110110    1001001010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37555 - 37559

  --1001001010111000    1001001010111001    1001001010111010    1001001010111011    1001001010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37560 - 37564

  --1001001010111101    1001001010111110    1001001010111111    1001001011000000    1001001011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37565 - 37569

  --1001001011000010    1001001011000011    1001001011000100    1001001011000101    1001001011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37570 - 37574

  --1001001011000111    1001001011001000    1001001011001001    1001001011001010    1001001011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37575 - 37579

  --1001001011001100    1001001011001101    1001001011001110    1001001011001111    1001001011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37580 - 37584

  --1001001011010001    1001001011010010    1001001011010011    1001001011010100    1001001011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37585 - 37589

  --1001001011010110    1001001011010111    1001001011011000    1001001011011001    1001001011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37590 - 37594

  --1001001011011011    1001001011011100    1001001011011101    1001001011011110    1001001011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37595 - 37599

  --1001001011100000    1001001011100001    1001001011100010    1001001011100011    1001001011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37600 - 37604

  --1001001011100101    1001001011100110    1001001011100111    1001001011101000    1001001011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37605 - 37609

  --1001001011101010    1001001011101011    1001001011101100    1001001011101101    1001001011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37610 - 37614

  --1001001011101111    1001001011110000    1001001011110001    1001001011110010    1001001011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37615 - 37619

  --1001001011110100    1001001011110101    1001001011110110    1001001011110111    1001001011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37620 - 37624

  --1001001011111001    1001001011111010    1001001011111011    1001001011111100    1001001011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37625 - 37629

  --1001001011111110    1001001011111111    1001001100000000    1001001100000001    1001001100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37630 - 37634

  --1001001100000011    1001001100000100    1001001100000101    1001001100000110    1001001100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37635 - 37639

  --1001001100001000    1001001100001001    1001001100001010    1001001100001011    1001001100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37640 - 37644

  --1001001100001101    1001001100001110    1001001100001111    1001001100010000    1001001100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37645 - 37649

  --1001001100010010    1001001100010011    1001001100010100    1001001100010101    1001001100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37650 - 37654

  --1001001100010111    1001001100011000    1001001100011001    1001001100011010    1001001100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37655 - 37659

  --1001001100011100    1001001100011101    1001001100011110    1001001100011111    1001001100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37660 - 37664

  --1001001100100001    1001001100100010    1001001100100011    1001001100100100    1001001100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37665 - 37669

  --1001001100100110    1001001100100111    1001001100101000    1001001100101001    1001001100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37670 - 37674

  --1001001100101011    1001001100101100    1001001100101101    1001001100101110    1001001100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37675 - 37679

  --1001001100110000    1001001100110001    1001001100110010    1001001100110011    1001001100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37680 - 37684

  --1001001100110101    1001001100110110    1001001100110111    1001001100111000    1001001100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37685 - 37689

  --1001001100111010    1001001100111011    1001001100111100    1001001100111101    1001001100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37690 - 37694

  --1001001100111111    1001001101000000    1001001101000001    1001001101000010    1001001101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37695 - 37699

  --1001001101000100    1001001101000101    1001001101000110    1001001101000111    1001001101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37700 - 37704

  --1001001101001001    1001001101001010    1001001101001011    1001001101001100    1001001101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37705 - 37709

  --1001001101001110    1001001101001111    1001001101010000    1001001101010001    1001001101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37710 - 37714

  --1001001101010011    1001001101010100    1001001101010101    1001001101010110    1001001101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37715 - 37719

  --1001001101011000    1001001101011001    1001001101011010    1001001101011011    1001001101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37720 - 37724

  --1001001101011101    1001001101011110    1001001101011111    1001001101100000    1001001101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37725 - 37729

  --1001001101100010    1001001101100011    1001001101100100    1001001101100101    1001001101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37730 - 37734

  --1001001101100111    1001001101101000    1001001101101001    1001001101101010    1001001101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37735 - 37739

  --1001001101101100    1001001101101101    1001001101101110    1001001101101111    1001001101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37740 - 37744

  --1001001101110001    1001001101110010    1001001101110011    1001001101110100    1001001101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37745 - 37749

  --1001001101110110    1001001101110111    1001001101111000    1001001101111001    1001001101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37750 - 37754

  --1001001101111011    1001001101111100    1001001101111101    1001001101111110    1001001101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37755 - 37759

  --1001001110000000    1001001110000001    1001001110000010    1001001110000011    1001001110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37760 - 37764

  --1001001110000101    1001001110000110    1001001110000111    1001001110001000    1001001110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37765 - 37769

  --1001001110001010    1001001110001011    1001001110001100    1001001110001101    1001001110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37770 - 37774

  --1001001110001111    1001001110010000    1001001110010001    1001001110010010    1001001110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37775 - 37779

  --1001001110010100    1001001110010101    1001001110010110    1001001110010111    1001001110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37780 - 37784

  --1001001110011001    1001001110011010    1001001110011011    1001001110011100    1001001110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37785 - 37789

  --1001001110011110    1001001110011111    1001001110100000    1001001110100001    1001001110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37790 - 37794

  --1001001110100011    1001001110100100    1001001110100101    1001001110100110    1001001110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37795 - 37799

  --1001001110101000    1001001110101001    1001001110101010    1001001110101011    1001001110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37800 - 37804

  --1001001110101101    1001001110101110    1001001110101111    1001001110110000    1001001110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37805 - 37809

  --1001001110110010    1001001110110011    1001001110110100    1001001110110101    1001001110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37810 - 37814

  --1001001110110111    1001001110111000    1001001110111001    1001001110111010    1001001110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37815 - 37819

  --1001001110111100    1001001110111101    1001001110111110    1001001110111111    1001001111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37820 - 37824

  --1001001111000001    1001001111000010    1001001111000011    1001001111000100    1001001111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37825 - 37829

  --1001001111000110    1001001111000111    1001001111001000    1001001111001001    1001001111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37830 - 37834

  --1001001111001011    1001001111001100    1001001111001101    1001001111001110    1001001111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37835 - 37839

  --1001001111010000    1001001111010001    1001001111010010    1001001111010011    1001001111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37840 - 37844

  --1001001111010101    1001001111010110    1001001111010111    1001001111011000    1001001111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37845 - 37849

  --1001001111011010    1001001111011011    1001001111011100    1001001111011101    1001001111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37850 - 37854

  --1001001111011111    1001001111100000    1001001111100001    1001001111100010    1001001111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37855 - 37859

  --1001001111100100    1001001111100101    1001001111100110    1001001111100111    1001001111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37860 - 37864

  --1001001111101001    1001001111101010    1001001111101011    1001001111101100    1001001111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37865 - 37869

  --1001001111101110    1001001111101111    1001001111110000    1001001111110001    1001001111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37870 - 37874

  --1001001111110011    1001001111110100    1001001111110101    1001001111110110    1001001111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37875 - 37879

  --1001001111111000    1001001111111001    1001001111111010    1001001111111011    1001001111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37880 - 37884

  --1001001111111101    1001001111111110    1001001111111111    1001010000000000    1001010000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37885 - 37889

  --1001010000000010    1001010000000011    1001010000000100    1001010000000101    1001010000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37890 - 37894

  --1001010000000111    1001010000001000    1001010000001001    1001010000001010    1001010000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37895 - 37899

  --1001010000001100    1001010000001101    1001010000001110    1001010000001111    1001010000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37900 - 37904

  --1001010000010001    1001010000010010    1001010000010011    1001010000010100    1001010000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37905 - 37909

  --1001010000010110    1001010000010111    1001010000011000    1001010000011001    1001010000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37910 - 37914

  --1001010000011011    1001010000011100    1001010000011101    1001010000011110    1001010000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37915 - 37919

  --1001010000100000    1001010000100001    1001010000100010    1001010000100011    1001010000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37920 - 37924

  --1001010000100101    1001010000100110    1001010000100111    1001010000101000    1001010000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37925 - 37929

  --1001010000101010    1001010000101011    1001010000101100    1001010000101101    1001010000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37930 - 37934

  --1001010000101111    1001010000110000    1001010000110001    1001010000110010    1001010000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37935 - 37939

  --1001010000110100    1001010000110101    1001010000110110    1001010000110111    1001010000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37940 - 37944

  --1001010000111001    1001010000111010    1001010000111011    1001010000111100    1001010000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37945 - 37949

  --1001010000111110    1001010000111111    1001010001000000    1001010001000001    1001010001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37950 - 37954

  --1001010001000011    1001010001000100    1001010001000101    1001010001000110    1001010001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37955 - 37959

  --1001010001001000    1001010001001001    1001010001001010    1001010001001011    1001010001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37960 - 37964

  --1001010001001101    1001010001001110    1001010001001111    1001010001010000    1001010001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37965 - 37969

  --1001010001010010    1001010001010011    1001010001010100    1001010001010101    1001010001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37970 - 37974

  --1001010001010111    1001010001011000    1001010001011001    1001010001011010    1001010001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37975 - 37979

  --1001010001011100    1001010001011101    1001010001011110    1001010001011111    1001010001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37980 - 37984

  --1001010001100001    1001010001100010    1001010001100011    1001010001100100    1001010001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37985 - 37989

  --1001010001100110    1001010001100111    1001010001101000    1001010001101001    1001010001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37990 - 37994

  --1001010001101011    1001010001101100    1001010001101101    1001010001101110    1001010001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 37995 - 37999

  --1001010001110000    1001010001110001    1001010001110010    1001010001110011    1001010001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38000 - 38004

  --1001010001110101    1001010001110110    1001010001110111    1001010001111000    1001010001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38005 - 38009

  --1001010001111010    1001010001111011    1001010001111100    1001010001111101    1001010001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38010 - 38014

  --1001010001111111    1001010010000000    1001010010000001    1001010010000010    1001010010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38015 - 38019

  --1001010010000100    1001010010000101    1001010010000110    1001010010000111    1001010010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38020 - 38024

  --1001010010001001    1001010010001010    1001010010001011    1001010010001100    1001010010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38025 - 38029

  --1001010010001110    1001010010001111    1001010010010000    1001010010010001    1001010010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38030 - 38034

  --1001010010010011    1001010010010100    1001010010010101    1001010010010110    1001010010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38035 - 38039

  --1001010010011000    1001010010011001    1001010010011010    1001010010011011    1001010010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38040 - 38044

  --1001010010011101    1001010010011110    1001010010011111    1001010010100000    1001010010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38045 - 38049

  --1001010010100010    1001010010100011    1001010010100100    1001010010100101    1001010010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38050 - 38054

  --1001010010100111    1001010010101000    1001010010101001    1001010010101010    1001010010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38055 - 38059

  --1001010010101100    1001010010101101    1001010010101110    1001010010101111    1001010010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38060 - 38064

  --1001010010110001    1001010010110010    1001010010110011    1001010010110100    1001010010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38065 - 38069

  --1001010010110110    1001010010110111    1001010010111000    1001010010111001    1001010010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38070 - 38074

  --1001010010111011    1001010010111100    1001010010111101    1001010010111110    1001010010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38075 - 38079

  --1001010011000000    1001010011000001    1001010011000010    1001010011000011    1001010011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38080 - 38084

  --1001010011000101    1001010011000110    1001010011000111    1001010011001000    1001010011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38085 - 38089

  --1001010011001010    1001010011001011    1001010011001100    1001010011001101    1001010011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38090 - 38094

  --1001010011001111    1001010011010000    1001010011010001    1001010011010010    1001010011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38095 - 38099

  --1001010011010100    1001010011010101    1001010011010110    1001010011010111    1001010011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38100 - 38104

  --1001010011011001    1001010011011010    1001010011011011    1001010011011100    1001010011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38105 - 38109

  --1001010011011110    1001010011011111    1001010011100000    1001010011100001    1001010011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38110 - 38114

  --1001010011100011    1001010011100100    1001010011100101    1001010011100110    1001010011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38115 - 38119

  --1001010011101000    1001010011101001    1001010011101010    1001010011101011    1001010011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38120 - 38124

  --1001010011101101    1001010011101110    1001010011101111    1001010011110000    1001010011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38125 - 38129

  --1001010011110010    1001010011110011    1001010011110100    1001010011110101    1001010011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38130 - 38134

  --1001010011110111    1001010011111000    1001010011111001    1001010011111010    1001010011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38135 - 38139

  --1001010011111100    1001010011111101    1001010011111110    1001010011111111    1001010100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38140 - 38144

  --1001010100000001    1001010100000010    1001010100000011    1001010100000100    1001010100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38145 - 38149

  --1001010100000110    1001010100000111    1001010100001000    1001010100001001    1001010100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38150 - 38154

  --1001010100001011    1001010100001100    1001010100001101    1001010100001110    1001010100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38155 - 38159

  --1001010100010000    1001010100010001    1001010100010010    1001010100010011    1001010100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38160 - 38164

  --1001010100010101    1001010100010110    1001010100010111    1001010100011000    1001010100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38165 - 38169

  --1001010100011010    1001010100011011    1001010100011100    1001010100011101    1001010100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38170 - 38174

  --1001010100011111    1001010100100000    1001010100100001    1001010100100010    1001010100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38175 - 38179

  --1001010100100100    1001010100100101    1001010100100110    1001010100100111    1001010100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38180 - 38184

  --1001010100101001    1001010100101010    1001010100101011    1001010100101100    1001010100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38185 - 38189

  --1001010100101110    1001010100101111    1001010100110000    1001010100110001    1001010100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38190 - 38194

  --1001010100110011    1001010100110100    1001010100110101    1001010100110110    1001010100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38195 - 38199

  --1001010100111000    1001010100111001    1001010100111010    1001010100111011    1001010100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38200 - 38204

  --1001010100111101    1001010100111110    1001010100111111    1001010101000000    1001010101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38205 - 38209

  --1001010101000010    1001010101000011    1001010101000100    1001010101000101    1001010101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38210 - 38214

  --1001010101000111    1001010101001000    1001010101001001    1001010101001010    1001010101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38215 - 38219

  --1001010101001100    1001010101001101    1001010101001110    1001010101001111    1001010101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38220 - 38224

  --1001010101010001    1001010101010010    1001010101010011    1001010101010100    1001010101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38225 - 38229

  --1001010101010110    1001010101010111    1001010101011000    1001010101011001    1001010101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38230 - 38234

  --1001010101011011    1001010101011100    1001010101011101    1001010101011110    1001010101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38235 - 38239

  --1001010101100000    1001010101100001    1001010101100010    1001010101100011    1001010101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38240 - 38244

  --1001010101100101    1001010101100110    1001010101100111    1001010101101000    1001010101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38245 - 38249

  --1001010101101010    1001010101101011    1001010101101100    1001010101101101    1001010101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38250 - 38254

  --1001010101101111    1001010101110000    1001010101110001    1001010101110010    1001010101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38255 - 38259

  --1001010101110100    1001010101110101    1001010101110110    1001010101110111    1001010101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38260 - 38264

  --1001010101111001    1001010101111010    1001010101111011    1001010101111100    1001010101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38265 - 38269

  --1001010101111110    1001010101111111    1001010110000000    1001010110000001    1001010110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38270 - 38274

  --1001010110000011    1001010110000100    1001010110000101    1001010110000110    1001010110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38275 - 38279

  --1001010110001000    1001010110001001    1001010110001010    1001010110001011    1001010110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38280 - 38284

  --1001010110001101    1001010110001110    1001010110001111    1001010110010000    1001010110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38285 - 38289

  --1001010110010010    1001010110010011    1001010110010100    1001010110010101    1001010110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38290 - 38294

  --1001010110010111    1001010110011000    1001010110011001    1001010110011010    1001010110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38295 - 38299

  --1001010110011100    1001010110011101    1001010110011110    1001010110011111    1001010110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38300 - 38304

  --1001010110100001    1001010110100010    1001010110100011    1001010110100100    1001010110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38305 - 38309

  --1001010110100110    1001010110100111    1001010110101000    1001010110101001    1001010110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38310 - 38314

  --1001010110101011    1001010110101100    1001010110101101    1001010110101110    1001010110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38315 - 38319

  --1001010110110000    1001010110110001    1001010110110010    1001010110110011    1001010110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38320 - 38324

  --1001010110110101    1001010110110110    1001010110110111    1001010110111000    1001010110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38325 - 38329

  --1001010110111010    1001010110111011    1001010110111100    1001010110111101    1001010110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38330 - 38334

  --1001010110111111    1001010111000000    1001010111000001    1001010111000010    1001010111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38335 - 38339

  --1001010111000100    1001010111000101    1001010111000110    1001010111000111    1001010111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38340 - 38344

  --1001010111001001    1001010111001010    1001010111001011    1001010111001100    1001010111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38345 - 38349

  --1001010111001110    1001010111001111    1001010111010000    1001010111010001    1001010111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38350 - 38354

  --1001010111010011    1001010111010100    1001010111010101    1001010111010110    1001010111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38355 - 38359

  --1001010111011000    1001010111011001    1001010111011010    1001010111011011    1001010111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38360 - 38364

  --1001010111011101    1001010111011110    1001010111011111    1001010111100000    1001010111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38365 - 38369

  --1001010111100010    1001010111100011    1001010111100100    1001010111100101    1001010111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38370 - 38374

  --1001010111100111    1001010111101000    1001010111101001    1001010111101010    1001010111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38375 - 38379

  --1001010111101100    1001010111101101    1001010111101110    1001010111101111    1001010111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38380 - 38384

  --1001010111110001    1001010111110010    1001010111110011    1001010111110100    1001010111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38385 - 38389

  --1001010111110110    1001010111110111    1001010111111000    1001010111111001    1001010111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38390 - 38394

  --1001010111111011    1001010111111100    1001010111111101    1001010111111110    1001010111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38395 - 38399

  --1001011000000000    1001011000000001    1001011000000010    1001011000000011    1001011000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38400 - 38404

  --1001011000000101    1001011000000110    1001011000000111    1001011000001000    1001011000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38405 - 38409

  --1001011000001010    1001011000001011    1001011000001100    1001011000001101    1001011000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38410 - 38414

  --1001011000001111    1001011000010000    1001011000010001    1001011000010010    1001011000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38415 - 38419

  --1001011000010100    1001011000010101    1001011000010110    1001011000010111    1001011000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38420 - 38424

  --1001011000011001    1001011000011010    1001011000011011    1001011000011100    1001011000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38425 - 38429

  --1001011000011110    1001011000011111    1001011000100000    1001011000100001    1001011000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38430 - 38434

  --1001011000100011    1001011000100100    1001011000100101    1001011000100110    1001011000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38435 - 38439

  --1001011000101000    1001011000101001    1001011000101010    1001011000101011    1001011000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38440 - 38444

  --1001011000101101    1001011000101110    1001011000101111    1001011000110000    1001011000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38445 - 38449

  --1001011000110010    1001011000110011    1001011000110100    1001011000110101    1001011000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38450 - 38454

  --1001011000110111    1001011000111000    1001011000111001    1001011000111010    1001011000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38455 - 38459

  --1001011000111100    1001011000111101    1001011000111110    1001011000111111    1001011001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38460 - 38464

  --1001011001000001    1001011001000010    1001011001000011    1001011001000100    1001011001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38465 - 38469

  --1001011001000110    1001011001000111    1001011001001000    1001011001001001    1001011001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38470 - 38474

  --1001011001001011    1001011001001100    1001011001001101    1001011001001110    1001011001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38475 - 38479

  --1001011001010000    1001011001010001    1001011001010010    1001011001010011    1001011001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38480 - 38484

  --1001011001010101    1001011001010110    1001011001010111    1001011001011000    1001011001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38485 - 38489

  --1001011001011010    1001011001011011    1001011001011100    1001011001011101    1001011001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38490 - 38494

  --1001011001011111    1001011001100000    1001011001100001    1001011001100010    1001011001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38495 - 38499

  --1001011001100100    1001011001100101    1001011001100110    1001011001100111    1001011001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38500 - 38504

  --1001011001101001    1001011001101010    1001011001101011    1001011001101100    1001011001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38505 - 38509

  --1001011001101110    1001011001101111    1001011001110000    1001011001110001    1001011001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38510 - 38514

  --1001011001110011    1001011001110100    1001011001110101    1001011001110110    1001011001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38515 - 38519

  --1001011001111000    1001011001111001    1001011001111010    1001011001111011    1001011001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38520 - 38524

  --1001011001111101    1001011001111110    1001011001111111    1001011010000000    1001011010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38525 - 38529

  --1001011010000010    1001011010000011    1001011010000100    1001011010000101    1001011010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38530 - 38534

  --1001011010000111    1001011010001000    1001011010001001    1001011010001010    1001011010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38535 - 38539

  --1001011010001100    1001011010001101    1001011010001110    1001011010001111    1001011010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38540 - 38544

  --1001011010010001    1001011010010010    1001011010010011    1001011010010100    1001011010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38545 - 38549

  --1001011010010110    1001011010010111    1001011010011000    1001011010011001    1001011010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38550 - 38554

  --1001011010011011    1001011010011100    1001011010011101    1001011010011110    1001011010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38555 - 38559

  --1001011010100000    1001011010100001    1001011010100010    1001011010100011    1001011010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38560 - 38564

  --1001011010100101    1001011010100110    1001011010100111    1001011010101000    1001011010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38565 - 38569

  --1001011010101010    1001011010101011    1001011010101100    1001011010101101    1001011010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38570 - 38574

  --1001011010101111    1001011010110000    1001011010110001    1001011010110010    1001011010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38575 - 38579

  --1001011010110100    1001011010110101    1001011010110110    1001011010110111    1001011010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38580 - 38584

  --1001011010111001    1001011010111010    1001011010111011    1001011010111100    1001011010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38585 - 38589

  --1001011010111110    1001011010111111    1001011011000000    1001011011000001    1001011011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38590 - 38594

  --1001011011000011    1001011011000100    1001011011000101    1001011011000110    1001011011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38595 - 38599

  --1001011011001000    1001011011001001    1001011011001010    1001011011001011    1001011011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38600 - 38604

  --1001011011001101    1001011011001110    1001011011001111    1001011011010000    1001011011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38605 - 38609

  --1001011011010010    1001011011010011    1001011011010100    1001011011010101    1001011011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38610 - 38614

  --1001011011010111    1001011011011000    1001011011011001    1001011011011010    1001011011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38615 - 38619

  --1001011011011100    1001011011011101    1001011011011110    1001011011011111    1001011011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38620 - 38624

  --1001011011100001    1001011011100010    1001011011100011    1001011011100100    1001011011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38625 - 38629

  --1001011011100110    1001011011100111    1001011011101000    1001011011101001    1001011011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38630 - 38634

  --1001011011101011    1001011011101100    1001011011101101    1001011011101110    1001011011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38635 - 38639

  --1001011011110000    1001011011110001    1001011011110010    1001011011110011    1001011011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38640 - 38644

  --1001011011110101    1001011011110110    1001011011110111    1001011011111000    1001011011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38645 - 38649

  --1001011011111010    1001011011111011    1001011011111100    1001011011111101    1001011011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38650 - 38654

  --1001011011111111    1001011100000000    1001011100000001    1001011100000010    1001011100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38655 - 38659

  --1001011100000100    1001011100000101    1001011100000110    1001011100000111    1001011100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38660 - 38664

  --1001011100001001    1001011100001010    1001011100001011    1001011100001100    1001011100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38665 - 38669

  --1001011100001110    1001011100001111    1001011100010000    1001011100010001    1001011100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38670 - 38674

  --1001011100010011    1001011100010100    1001011100010101    1001011100010110    1001011100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38675 - 38679

  --1001011100011000    1001011100011001    1001011100011010    1001011100011011    1001011100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38680 - 38684

  --1001011100011101    1001011100011110    1001011100011111    1001011100100000    1001011100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38685 - 38689

  --1001011100100010    1001011100100011    1001011100100100    1001011100100101    1001011100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38690 - 38694

  --1001011100100111    1001011100101000    1001011100101001    1001011100101010    1001011100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38695 - 38699

  --1001011100101100    1001011100101101    1001011100101110    1001011100101111    1001011100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38700 - 38704

  --1001011100110001    1001011100110010    1001011100110011    1001011100110100    1001011100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38705 - 38709

  --1001011100110110    1001011100110111    1001011100111000    1001011100111001    1001011100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38710 - 38714

  --1001011100111011    1001011100111100    1001011100111101    1001011100111110    1001011100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38715 - 38719

  --1001011101000000    1001011101000001    1001011101000010    1001011101000011    1001011101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38720 - 38724

  --1001011101000101    1001011101000110    1001011101000111    1001011101001000    1001011101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38725 - 38729

  --1001011101001010    1001011101001011    1001011101001100    1001011101001101    1001011101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38730 - 38734

  --1001011101001111    1001011101010000    1001011101010001    1001011101010010    1001011101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38735 - 38739

  --1001011101010100    1001011101010101    1001011101010110    1001011101010111    1001011101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38740 - 38744

  --1001011101011001    1001011101011010    1001011101011011    1001011101011100    1001011101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38745 - 38749

  --1001011101011110    1001011101011111    1001011101100000    1001011101100001    1001011101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38750 - 38754

  --1001011101100011    1001011101100100    1001011101100101    1001011101100110    1001011101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38755 - 38759

  --1001011101101000    1001011101101001    1001011101101010    1001011101101011    1001011101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38760 - 38764

  --1001011101101101    1001011101101110    1001011101101111    1001011101110000    1001011101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38765 - 38769

  --1001011101110010    1001011101110011    1001011101110100    1001011101110101    1001011101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38770 - 38774

  --1001011101110111    1001011101111000    1001011101111001    1001011101111010    1001011101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38775 - 38779

  --1001011101111100    1001011101111101    1001011101111110    1001011101111111    1001011110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38780 - 38784

  --1001011110000001    1001011110000010    1001011110000011    1001011110000100    1001011110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38785 - 38789

  --1001011110000110    1001011110000111    1001011110001000    1001011110001001    1001011110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38790 - 38794

  --1001011110001011    1001011110001100    1001011110001101    1001011110001110    1001011110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38795 - 38799

  --1001011110010000    1001011110010001    1001011110010010    1001011110010011    1001011110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38800 - 38804

  --1001011110010101    1001011110010110    1001011110010111    1001011110011000    1001011110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38805 - 38809

  --1001011110011010    1001011110011011    1001011110011100    1001011110011101    1001011110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38810 - 38814

  --1001011110011111    1001011110100000    1001011110100001    1001011110100010    1001011110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38815 - 38819

  --1001011110100100    1001011110100101    1001011110100110    1001011110100111    1001011110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38820 - 38824

  --1001011110101001    1001011110101010    1001011110101011    1001011110101100    1001011110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38825 - 38829

  --1001011110101110    1001011110101111    1001011110110000    1001011110110001    1001011110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38830 - 38834

  --1001011110110011    1001011110110100    1001011110110101    1001011110110110    1001011110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38835 - 38839

  --1001011110111000    1001011110111001    1001011110111010    1001011110111011    1001011110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38840 - 38844

  --1001011110111101    1001011110111110    1001011110111111    1001011111000000    1001011111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38845 - 38849

  --1001011111000010    1001011111000011    1001011111000100    1001011111000101    1001011111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38850 - 38854

  --1001011111000111    1001011111001000    1001011111001001    1001011111001010    1001011111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38855 - 38859

  --1001011111001100    1001011111001101    1001011111001110    1001011111001111    1001011111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38860 - 38864

  --1001011111010001    1001011111010010    1001011111010011    1001011111010100    1001011111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38865 - 38869

  --1001011111010110    1001011111010111    1001011111011000    1001011111011001    1001011111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38870 - 38874

  --1001011111011011    1001011111011100    1001011111011101    1001011111011110    1001011111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38875 - 38879

  --1001011111100000    1001011111100001    1001011111100010    1001011111100011    1001011111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38880 - 38884

  --1001011111100101    1001011111100110    1001011111100111    1001011111101000    1001011111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38885 - 38889

  --1001011111101010    1001011111101011    1001011111101100    1001011111101101    1001011111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38890 - 38894

  --1001011111101111    1001011111110000    1001011111110001    1001011111110010    1001011111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38895 - 38899

  --1001011111110100    1001011111110101    1001011111110110    1001011111110111    1001011111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38900 - 38904

  --1001011111111001    1001011111111010    1001011111111011    1001011111111100    1001011111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38905 - 38909

  --1001011111111110    1001011111111111    1001100000000000    1001100000000001    1001100000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38910 - 38914

  --1001100000000011    1001100000000100    1001100000000101    1001100000000110    1001100000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38915 - 38919

  --1001100000001000    1001100000001001    1001100000001010    1001100000001011    1001100000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38920 - 38924

  --1001100000001101    1001100000001110    1001100000001111    1001100000010000    1001100000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38925 - 38929

  --1001100000010010    1001100000010011    1001100000010100    1001100000010101    1001100000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38930 - 38934

  --1001100000010111    1001100000011000    1001100000011001    1001100000011010    1001100000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38935 - 38939

  --1001100000011100    1001100000011101    1001100000011110    1001100000011111    1001100000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38940 - 38944

  --1001100000100001    1001100000100010    1001100000100011    1001100000100100    1001100000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38945 - 38949

  --1001100000100110    1001100000100111    1001100000101000    1001100000101001    1001100000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38950 - 38954

  --1001100000101011    1001100000101100    1001100000101101    1001100000101110    1001100000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38955 - 38959

  --1001100000110000    1001100000110001    1001100000110010    1001100000110011    1001100000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38960 - 38964

  --1001100000110101    1001100000110110    1001100000110111    1001100000111000    1001100000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38965 - 38969

  --1001100000111010    1001100000111011    1001100000111100    1001100000111101    1001100000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38970 - 38974

  --1001100000111111    1001100001000000    1001100001000001    1001100001000010    1001100001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38975 - 38979

  --1001100001000100    1001100001000101    1001100001000110    1001100001000111    1001100001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38980 - 38984

  --1001100001001001    1001100001001010    1001100001001011    1001100001001100    1001100001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38985 - 38989

  --1001100001001110    1001100001001111    1001100001010000    1001100001010001    1001100001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38990 - 38994

  --1001100001010011    1001100001010100    1001100001010101    1001100001010110    1001100001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 38995 - 38999

  --1001100001011000    1001100001011001    1001100001011010    1001100001011011    1001100001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39000 - 39004

  --1001100001011101    1001100001011110    1001100001011111    1001100001100000    1001100001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39005 - 39009

  --1001100001100010    1001100001100011    1001100001100100    1001100001100101    1001100001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39010 - 39014

  --1001100001100111    1001100001101000    1001100001101001    1001100001101010    1001100001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39015 - 39019

  --1001100001101100    1001100001101101    1001100001101110    1001100001101111    1001100001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39020 - 39024

  --1001100001110001    1001100001110010    1001100001110011    1001100001110100    1001100001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39025 - 39029

  --1001100001110110    1001100001110111    1001100001111000    1001100001111001    1001100001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39030 - 39034

  --1001100001111011    1001100001111100    1001100001111101    1001100001111110    1001100001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39035 - 39039

  --1001100010000000    1001100010000001    1001100010000010    1001100010000011    1001100010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39040 - 39044

  --1001100010000101    1001100010000110    1001100010000111    1001100010001000    1001100010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39045 - 39049

  --1001100010001010    1001100010001011    1001100010001100    1001100010001101    1001100010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39050 - 39054

  --1001100010001111    1001100010010000    1001100010010001    1001100010010010    1001100010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39055 - 39059

  --1001100010010100    1001100010010101    1001100010010110    1001100010010111    1001100010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39060 - 39064

  --1001100010011001    1001100010011010    1001100010011011    1001100010011100    1001100010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39065 - 39069

  --1001100010011110    1001100010011111    1001100010100000    1001100010100001    1001100010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39070 - 39074

  --1001100010100011    1001100010100100    1001100010100101    1001100010100110    1001100010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39075 - 39079

  --1001100010101000    1001100010101001    1001100010101010    1001100010101011    1001100010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39080 - 39084

  --1001100010101101    1001100010101110    1001100010101111    1001100010110000    1001100010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39085 - 39089

  --1001100010110010    1001100010110011    1001100010110100    1001100010110101    1001100010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39090 - 39094

  --1001100010110111    1001100010111000    1001100010111001    1001100010111010    1001100010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39095 - 39099

  --1001100010111100    1001100010111101    1001100010111110    1001100010111111    1001100011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39100 - 39104

  --1001100011000001    1001100011000010    1001100011000011    1001100011000100    1001100011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39105 - 39109

  --1001100011000110    1001100011000111    1001100011001000    1001100011001001    1001100011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39110 - 39114

  --1001100011001011    1001100011001100    1001100011001101    1001100011001110    1001100011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39115 - 39119

  --1001100011010000    1001100011010001    1001100011010010    1001100011010011    1001100011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39120 - 39124

  --1001100011010101    1001100011010110    1001100011010111    1001100011011000    1001100011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39125 - 39129

  --1001100011011010    1001100011011011    1001100011011100    1001100011011101    1001100011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39130 - 39134

  --1001100011011111    1001100011100000    1001100011100001    1001100011100010    1001100011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39135 - 39139

  --1001100011100100    1001100011100101    1001100011100110    1001100011100111    1001100011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39140 - 39144

  --1001100011101001    1001100011101010    1001100011101011    1001100011101100    1001100011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39145 - 39149

  --1001100011101110    1001100011101111    1001100011110000    1001100011110001    1001100011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39150 - 39154

  --1001100011110011    1001100011110100    1001100011110101    1001100011110110    1001100011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39155 - 39159

  --1001100011111000    1001100011111001    1001100011111010    1001100011111011    1001100011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39160 - 39164

  --1001100011111101    1001100011111110    1001100011111111    1001100100000000    1001100100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39165 - 39169

  --1001100100000010    1001100100000011    1001100100000100    1001100100000101    1001100100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39170 - 39174

  --1001100100000111    1001100100001000    1001100100001001    1001100100001010    1001100100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39175 - 39179

  --1001100100001100    1001100100001101    1001100100001110    1001100100001111    1001100100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39180 - 39184

  --1001100100010001    1001100100010010    1001100100010011    1001100100010100    1001100100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39185 - 39189

  --1001100100010110    1001100100010111    1001100100011000    1001100100011001    1001100100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39190 - 39194

  --1001100100011011    1001100100011100    1001100100011101    1001100100011110    1001100100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39195 - 39199

  --1001100100100000    1001100100100001    1001100100100010    1001100100100011    1001100100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39200 - 39204

  --1001100100100101    1001100100100110    1001100100100111    1001100100101000    1001100100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39205 - 39209

  --1001100100101010    1001100100101011    1001100100101100    1001100100101101    1001100100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39210 - 39214

  --1001100100101111    1001100100110000    1001100100110001    1001100100110010    1001100100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39215 - 39219

  --1001100100110100    1001100100110101    1001100100110110    1001100100110111    1001100100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39220 - 39224

  --1001100100111001    1001100100111010    1001100100111011    1001100100111100    1001100100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39225 - 39229

  --1001100100111110    1001100100111111    1001100101000000    1001100101000001    1001100101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39230 - 39234

  --1001100101000011    1001100101000100    1001100101000101    1001100101000110    1001100101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39235 - 39239

  --1001100101001000    1001100101001001    1001100101001010    1001100101001011    1001100101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39240 - 39244

  --1001100101001101    1001100101001110    1001100101001111    1001100101010000    1001100101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39245 - 39249

  --1001100101010010    1001100101010011    1001100101010100    1001100101010101    1001100101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39250 - 39254

  --1001100101010111    1001100101011000    1001100101011001    1001100101011010    1001100101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39255 - 39259

  --1001100101011100    1001100101011101    1001100101011110    1001100101011111    1001100101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39260 - 39264

  --1001100101100001    1001100101100010    1001100101100011    1001100101100100    1001100101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39265 - 39269

  --1001100101100110    1001100101100111    1001100101101000    1001100101101001    1001100101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39270 - 39274

  --1001100101101011    1001100101101100    1001100101101101    1001100101101110    1001100101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39275 - 39279

  --1001100101110000    1001100101110001    1001100101110010    1001100101110011    1001100101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39280 - 39284

  --1001100101110101    1001100101110110    1001100101110111    1001100101111000    1001100101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39285 - 39289

  --1001100101111010    1001100101111011    1001100101111100    1001100101111101    1001100101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39290 - 39294

  --1001100101111111    1001100110000000    1001100110000001    1001100110000010    1001100110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39295 - 39299

  --1001100110000100    1001100110000101    1001100110000110    1001100110000111    1001100110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39300 - 39304

  --1001100110001001    1001100110001010    1001100110001011    1001100110001100    1001100110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39305 - 39309

  --1001100110001110    1001100110001111    1001100110010000    1001100110010001    1001100110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39310 - 39314

  --1001100110010011    1001100110010100    1001100110010101    1001100110010110    1001100110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39315 - 39319

  --1001100110011000    1001100110011001    1001100110011010    1001100110011011    1001100110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39320 - 39324

  --1001100110011101    1001100110011110    1001100110011111    1001100110100000    1001100110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39325 - 39329

  --1001100110100010    1001100110100011    1001100110100100    1001100110100101    1001100110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39330 - 39334

  --1001100110100111    1001100110101000    1001100110101001    1001100110101010    1001100110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39335 - 39339

  --1001100110101100    1001100110101101    1001100110101110    1001100110101111    1001100110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39340 - 39344

  --1001100110110001    1001100110110010    1001100110110011    1001100110110100    1001100110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39345 - 39349

  --1001100110110110    1001100110110111    1001100110111000    1001100110111001    1001100110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39350 - 39354

  --1001100110111011    1001100110111100    1001100110111101    1001100110111110    1001100110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39355 - 39359

  --1001100111000000    1001100111000001    1001100111000010    1001100111000011    1001100111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39360 - 39364

  --1001100111000101    1001100111000110    1001100111000111    1001100111001000    1001100111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39365 - 39369

  --1001100111001010    1001100111001011    1001100111001100    1001100111001101    1001100111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39370 - 39374

  --1001100111001111    1001100111010000    1001100111010001    1001100111010010    1001100111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39375 - 39379

  --1001100111010100    1001100111010101    1001100111010110    1001100111010111    1001100111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39380 - 39384

  --1001100111011001    1001100111011010    1001100111011011    1001100111011100    1001100111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39385 - 39389

  --1001100111011110    1001100111011111    1001100111100000    1001100111100001    1001100111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39390 - 39394

  --1001100111100011    1001100111100100    1001100111100101    1001100111100110    1001100111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39395 - 39399

  --1001100111101000    1001100111101001    1001100111101010    1001100111101011    1001100111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39400 - 39404

  --1001100111101101    1001100111101110    1001100111101111    1001100111110000    1001100111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39405 - 39409

  --1001100111110010    1001100111110011    1001100111110100    1001100111110101    1001100111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39410 - 39414

  --1001100111110111    1001100111111000    1001100111111001    1001100111111010    1001100111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39415 - 39419

  --1001100111111100    1001100111111101    1001100111111110    1001100111111111    1001101000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39420 - 39424

  --1001101000000001    1001101000000010    1001101000000011    1001101000000100    1001101000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39425 - 39429

  --1001101000000110    1001101000000111    1001101000001000    1001101000001001    1001101000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39430 - 39434

  --1001101000001011    1001101000001100    1001101000001101    1001101000001110    1001101000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39435 - 39439

  --1001101000010000    1001101000010001    1001101000010010    1001101000010011    1001101000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39440 - 39444

  --1001101000010101    1001101000010110    1001101000010111    1001101000011000    1001101000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39445 - 39449

  --1001101000011010    1001101000011011    1001101000011100    1001101000011101    1001101000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39450 - 39454

  --1001101000011111    1001101000100000    1001101000100001    1001101000100010    1001101000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39455 - 39459

  --1001101000100100    1001101000100101    1001101000100110    1001101000100111    1001101000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39460 - 39464

  --1001101000101001    1001101000101010    1001101000101011    1001101000101100    1001101000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39465 - 39469

  --1001101000101110    1001101000101111    1001101000110000    1001101000110001    1001101000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39470 - 39474

  --1001101000110011    1001101000110100    1001101000110101    1001101000110110    1001101000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39475 - 39479

  --1001101000111000    1001101000111001    1001101000111010    1001101000111011    1001101000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39480 - 39484

  --1001101000111101    1001101000111110    1001101000111111    1001101001000000    1001101001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39485 - 39489

  --1001101001000010    1001101001000011    1001101001000100    1001101001000101    1001101001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39490 - 39494

  --1001101001000111    1001101001001000    1001101001001001    1001101001001010    1001101001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39495 - 39499

  --1001101001001100    1001101001001101    1001101001001110    1001101001001111    1001101001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39500 - 39504

  --1001101001010001    1001101001010010    1001101001010011    1001101001010100    1001101001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39505 - 39509

  --1001101001010110    1001101001010111    1001101001011000    1001101001011001    1001101001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39510 - 39514

  --1001101001011011    1001101001011100    1001101001011101    1001101001011110    1001101001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39515 - 39519

  --1001101001100000    1001101001100001    1001101001100010    1001101001100011    1001101001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39520 - 39524

  --1001101001100101    1001101001100110    1001101001100111    1001101001101000    1001101001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39525 - 39529

  --1001101001101010    1001101001101011    1001101001101100    1001101001101101    1001101001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39530 - 39534

  --1001101001101111    1001101001110000    1001101001110001    1001101001110010    1001101001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39535 - 39539

  --1001101001110100    1001101001110101    1001101001110110    1001101001110111    1001101001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39540 - 39544

  --1001101001111001    1001101001111010    1001101001111011    1001101001111100    1001101001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39545 - 39549

  --1001101001111110    1001101001111111    1001101010000000    1001101010000001    1001101010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39550 - 39554

  --1001101010000011    1001101010000100    1001101010000101    1001101010000110    1001101010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39555 - 39559

  --1001101010001000    1001101010001001    1001101010001010    1001101010001011    1001101010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39560 - 39564

  --1001101010001101    1001101010001110    1001101010001111    1001101010010000    1001101010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39565 - 39569

  --1001101010010010    1001101010010011    1001101010010100    1001101010010101    1001101010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39570 - 39574

  --1001101010010111    1001101010011000    1001101010011001    1001101010011010    1001101010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39575 - 39579

  --1001101010011100    1001101010011101    1001101010011110    1001101010011111    1001101010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39580 - 39584

  --1001101010100001    1001101010100010    1001101010100011    1001101010100100    1001101010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39585 - 39589

  --1001101010100110    1001101010100111    1001101010101000    1001101010101001    1001101010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39590 - 39594

  --1001101010101011    1001101010101100    1001101010101101    1001101010101110    1001101010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39595 - 39599

  --1001101010110000    1001101010110001    1001101010110010    1001101010110011    1001101010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39600 - 39604

  --1001101010110101    1001101010110110    1001101010110111    1001101010111000    1001101010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39605 - 39609

  --1001101010111010    1001101010111011    1001101010111100    1001101010111101    1001101010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39610 - 39614

  --1001101010111111    1001101011000000    1001101011000001    1001101011000010    1001101011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39615 - 39619

  --1001101011000100    1001101011000101    1001101011000110    1001101011000111    1001101011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39620 - 39624

  --1001101011001001    1001101011001010    1001101011001011    1001101011001100    1001101011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39625 - 39629

  --1001101011001110    1001101011001111    1001101011010000    1001101011010001    1001101011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39630 - 39634

  --1001101011010011    1001101011010100    1001101011010101    1001101011010110    1001101011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39635 - 39639

  --1001101011011000    1001101011011001    1001101011011010    1001101011011011    1001101011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39640 - 39644

  --1001101011011101    1001101011011110    1001101011011111    1001101011100000    1001101011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39645 - 39649

  --1001101011100010    1001101011100011    1001101011100100    1001101011100101    1001101011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39650 - 39654

  --1001101011100111    1001101011101000    1001101011101001    1001101011101010    1001101011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39655 - 39659

  --1001101011101100    1001101011101101    1001101011101110    1001101011101111    1001101011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39660 - 39664

  --1001101011110001    1001101011110010    1001101011110011    1001101011110100    1001101011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39665 - 39669

  --1001101011110110    1001101011110111    1001101011111000    1001101011111001    1001101011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39670 - 39674

  --1001101011111011    1001101011111100    1001101011111101    1001101011111110    1001101011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39675 - 39679

  --1001101100000000    1001101100000001    1001101100000010    1001101100000011    1001101100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39680 - 39684

  --1001101100000101    1001101100000110    1001101100000111    1001101100001000    1001101100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39685 - 39689

  --1001101100001010    1001101100001011    1001101100001100    1001101100001101    1001101100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39690 - 39694

  --1001101100001111    1001101100010000    1001101100010001    1001101100010010    1001101100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39695 - 39699

  --1001101100010100    1001101100010101    1001101100010110    1001101100010111    1001101100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39700 - 39704

  --1001101100011001    1001101100011010    1001101100011011    1001101100011100    1001101100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39705 - 39709

  --1001101100011110    1001101100011111    1001101100100000    1001101100100001    1001101100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39710 - 39714

  --1001101100100011    1001101100100100    1001101100100101    1001101100100110    1001101100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39715 - 39719

  --1001101100101000    1001101100101001    1001101100101010    1001101100101011    1001101100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39720 - 39724

  --1001101100101101    1001101100101110    1001101100101111    1001101100110000    1001101100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39725 - 39729

  --1001101100110010    1001101100110011    1001101100110100    1001101100110101    1001101100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39730 - 39734

  --1001101100110111    1001101100111000    1001101100111001    1001101100111010    1001101100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39735 - 39739

  --1001101100111100    1001101100111101    1001101100111110    1001101100111111    1001101101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39740 - 39744

  --1001101101000001    1001101101000010    1001101101000011    1001101101000100    1001101101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39745 - 39749

  --1001101101000110    1001101101000111    1001101101001000    1001101101001001    1001101101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39750 - 39754

  --1001101101001011    1001101101001100    1001101101001101    1001101101001110    1001101101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39755 - 39759

  --1001101101010000    1001101101010001    1001101101010010    1001101101010011    1001101101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39760 - 39764

  --1001101101010101    1001101101010110    1001101101010111    1001101101011000    1001101101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39765 - 39769

  --1001101101011010    1001101101011011    1001101101011100    1001101101011101    1001101101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39770 - 39774

  --1001101101011111    1001101101100000    1001101101100001    1001101101100010    1001101101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39775 - 39779

  --1001101101100100    1001101101100101    1001101101100110    1001101101100111    1001101101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39780 - 39784

  --1001101101101001    1001101101101010    1001101101101011    1001101101101100    1001101101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39785 - 39789

  --1001101101101110    1001101101101111    1001101101110000    1001101101110001    1001101101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39790 - 39794

  --1001101101110011    1001101101110100    1001101101110101    1001101101110110    1001101101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39795 - 39799

  --1001101101111000    1001101101111001    1001101101111010    1001101101111011    1001101101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39800 - 39804

  --1001101101111101    1001101101111110    1001101101111111    1001101110000000    1001101110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39805 - 39809

  --1001101110000010    1001101110000011    1001101110000100    1001101110000101    1001101110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39810 - 39814

  --1001101110000111    1001101110001000    1001101110001001    1001101110001010    1001101110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39815 - 39819

  --1001101110001100    1001101110001101    1001101110001110    1001101110001111    1001101110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39820 - 39824

  --1001101110010001    1001101110010010    1001101110010011    1001101110010100    1001101110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39825 - 39829

  --1001101110010110    1001101110010111    1001101110011000    1001101110011001    1001101110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39830 - 39834

  --1001101110011011    1001101110011100    1001101110011101    1001101110011110    1001101110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39835 - 39839

  --1001101110100000    1001101110100001    1001101110100010    1001101110100011    1001101110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39840 - 39844

  --1001101110100101    1001101110100110    1001101110100111    1001101110101000    1001101110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39845 - 39849

  --1001101110101010    1001101110101011    1001101110101100    1001101110101101    1001101110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39850 - 39854

  --1001101110101111    1001101110110000    1001101110110001    1001101110110010    1001101110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39855 - 39859

  --1001101110110100    1001101110110101    1001101110110110    1001101110110111    1001101110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39860 - 39864

  --1001101110111001    1001101110111010    1001101110111011    1001101110111100    1001101110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39865 - 39869

  --1001101110111110    1001101110111111    1001101111000000    1001101111000001    1001101111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39870 - 39874

  --1001101111000011    1001101111000100    1001101111000101    1001101111000110    1001101111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39875 - 39879

  --1001101111001000    1001101111001001    1001101111001010    1001101111001011    1001101111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39880 - 39884

  --1001101111001101    1001101111001110    1001101111001111    1001101111010000    1001101111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39885 - 39889

  --1001101111010010    1001101111010011    1001101111010100    1001101111010101    1001101111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39890 - 39894

  --1001101111010111    1001101111011000    1001101111011001    1001101111011010    1001101111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39895 - 39899

  --1001101111011100    1001101111011101    1001101111011110    1001101111011111    1001101111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39900 - 39904

  --1001101111100001    1001101111100010    1001101111100011    1001101111100100    1001101111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39905 - 39909

  --1001101111100110    1001101111100111    1001101111101000    1001101111101001    1001101111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39910 - 39914

  --1001101111101011    1001101111101100    1001101111101101    1001101111101110    1001101111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39915 - 39919

  --1001101111110000    1001101111110001    1001101111110010    1001101111110011    1001101111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39920 - 39924

  --1001101111110101    1001101111110110    1001101111110111    1001101111111000    1001101111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39925 - 39929

  --1001101111111010    1001101111111011    1001101111111100    1001101111111101    1001101111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39930 - 39934

  --1001101111111111    1001110000000000    1001110000000001    1001110000000010    1001110000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39935 - 39939

  --1001110000000100    1001110000000101    1001110000000110    1001110000000111    1001110000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39940 - 39944

  --1001110000001001    1001110000001010    1001110000001011    1001110000001100    1001110000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39945 - 39949

  --1001110000001110    1001110000001111    1001110000010000    1001110000010001    1001110000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39950 - 39954

  --1001110000010011    1001110000010100    1001110000010101    1001110000010110    1001110000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39955 - 39959

  --1001110000011000    1001110000011001    1001110000011010    1001110000011011    1001110000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39960 - 39964

  --1001110000011101    1001110000011110    1001110000011111    1001110000100000    1001110000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39965 - 39969

  --1001110000100010    1001110000100011    1001110000100100    1001110000100101    1001110000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39970 - 39974

  --1001110000100111    1001110000101000    1001110000101001    1001110000101010    1001110000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39975 - 39979

  --1001110000101100    1001110000101101    1001110000101110    1001110000101111    1001110000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39980 - 39984

  --1001110000110001    1001110000110010    1001110000110011    1001110000110100    1001110000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39985 - 39989

  --1001110000110110    1001110000110111    1001110000111000    1001110000111001    1001110000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39990 - 39994

  --1001110000111011    1001110000111100    1001110000111101    1001110000111110    1001110000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 39995 - 39999

  --1001110001000000    1001110001000001    1001110001000010    1001110001000011    1001110001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40000 - 40004

  --1001110001000101    1001110001000110    1001110001000111    1001110001001000    1001110001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40005 - 40009

  --1001110001001010    1001110001001011    1001110001001100    1001110001001101    1001110001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40010 - 40014

  --1001110001001111    1001110001010000    1001110001010001    1001110001010010    1001110001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40015 - 40019

  --1001110001010100    1001110001010101    1001110001010110    1001110001010111    1001110001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40020 - 40024

  --1001110001011001    1001110001011010    1001110001011011    1001110001011100    1001110001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40025 - 40029

  --1001110001011110    1001110001011111    1001110001100000    1001110001100001    1001110001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40030 - 40034

  --1001110001100011    1001110001100100    1001110001100101    1001110001100110    1001110001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40035 - 40039

  --1001110001101000    1001110001101001    1001110001101010    1001110001101011    1001110001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40040 - 40044

  --1001110001101101    1001110001101110    1001110001101111    1001110001110000    1001110001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40045 - 40049

  --1001110001110010    1001110001110011    1001110001110100    1001110001110101    1001110001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40050 - 40054

  --1001110001110111    1001110001111000    1001110001111001    1001110001111010    1001110001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40055 - 40059

  --1001110001111100    1001110001111101    1001110001111110    1001110001111111    1001110010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40060 - 40064

  --1001110010000001    1001110010000010    1001110010000011    1001110010000100    1001110010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40065 - 40069

  --1001110010000110    1001110010000111    1001110010001000    1001110010001001    1001110010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40070 - 40074

  --1001110010001011    1001110010001100    1001110010001101    1001110010001110    1001110010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40075 - 40079

  --1001110010010000    1001110010010001    1001110010010010    1001110010010011    1001110010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40080 - 40084

  --1001110010010101    1001110010010110    1001110010010111    1001110010011000    1001110010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40085 - 40089

  --1001110010011010    1001110010011011    1001110010011100    1001110010011101    1001110010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40090 - 40094

  --1001110010011111    1001110010100000    1001110010100001    1001110010100010    1001110010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40095 - 40099

  --1001110010100100    1001110010100101    1001110010100110    1001110010100111    1001110010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40100 - 40104

  --1001110010101001    1001110010101010    1001110010101011    1001110010101100    1001110010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40105 - 40109

  --1001110010101110    1001110010101111    1001110010110000    1001110010110001    1001110010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40110 - 40114

  --1001110010110011    1001110010110100    1001110010110101    1001110010110110    1001110010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40115 - 40119

  --1001110010111000    1001110010111001    1001110010111010    1001110010111011    1001110010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40120 - 40124

  --1001110010111101    1001110010111110    1001110010111111    1001110011000000    1001110011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40125 - 40129

  --1001110011000010    1001110011000011    1001110011000100    1001110011000101    1001110011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40130 - 40134

  --1001110011000111    1001110011001000    1001110011001001    1001110011001010    1001110011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40135 - 40139

  --1001110011001100    1001110011001101    1001110011001110    1001110011001111    1001110011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40140 - 40144

  --1001110011010001    1001110011010010    1001110011010011    1001110011010100    1001110011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40145 - 40149

  --1001110011010110    1001110011010111    1001110011011000    1001110011011001    1001110011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40150 - 40154

  --1001110011011011    1001110011011100    1001110011011101    1001110011011110    1001110011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40155 - 40159

  --1001110011100000    1001110011100001    1001110011100010    1001110011100011    1001110011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40160 - 40164

  --1001110011100101    1001110011100110    1001110011100111    1001110011101000    1001110011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40165 - 40169

  --1001110011101010    1001110011101011    1001110011101100    1001110011101101    1001110011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40170 - 40174

  --1001110011101111    1001110011110000    1001110011110001    1001110011110010    1001110011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40175 - 40179

  --1001110011110100    1001110011110101    1001110011110110    1001110011110111    1001110011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40180 - 40184

  --1001110011111001    1001110011111010    1001110011111011    1001110011111100    1001110011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40185 - 40189

  --1001110011111110    1001110011111111    1001110100000000    1001110100000001    1001110100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40190 - 40194

  --1001110100000011    1001110100000100    1001110100000101    1001110100000110    1001110100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40195 - 40199

  --1001110100001000    1001110100001001    1001110100001010    1001110100001011    1001110100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40200 - 40204

  --1001110100001101    1001110100001110    1001110100001111    1001110100010000    1001110100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40205 - 40209

  --1001110100010010    1001110100010011    1001110100010100    1001110100010101    1001110100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40210 - 40214

  --1001110100010111    1001110100011000    1001110100011001    1001110100011010    1001110100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40215 - 40219

  --1001110100011100    1001110100011101    1001110100011110    1001110100011111    1001110100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40220 - 40224

  --1001110100100001    1001110100100010    1001110100100011    1001110100100100    1001110100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40225 - 40229

  --1001110100100110    1001110100100111    1001110100101000    1001110100101001    1001110100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40230 - 40234

  --1001110100101011    1001110100101100    1001110100101101    1001110100101110    1001110100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40235 - 40239

  --1001110100110000    1001110100110001    1001110100110010    1001110100110011    1001110100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40240 - 40244

  --1001110100110101    1001110100110110    1001110100110111    1001110100111000    1001110100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40245 - 40249

  --1001110100111010    1001110100111011    1001110100111100    1001110100111101    1001110100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40250 - 40254

  --1001110100111111    1001110101000000    1001110101000001    1001110101000010    1001110101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40255 - 40259

  --1001110101000100    1001110101000101    1001110101000110    1001110101000111    1001110101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40260 - 40264

  --1001110101001001    1001110101001010    1001110101001011    1001110101001100    1001110101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40265 - 40269

  --1001110101001110    1001110101001111    1001110101010000    1001110101010001    1001110101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40270 - 40274

  --1001110101010011    1001110101010100    1001110101010101    1001110101010110    1001110101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40275 - 40279

  --1001110101011000    1001110101011001    1001110101011010    1001110101011011    1001110101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40280 - 40284

  --1001110101011101    1001110101011110    1001110101011111    1001110101100000    1001110101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40285 - 40289

  --1001110101100010    1001110101100011    1001110101100100    1001110101100101    1001110101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40290 - 40294

  --1001110101100111    1001110101101000    1001110101101001    1001110101101010    1001110101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40295 - 40299

  --1001110101101100    1001110101101101    1001110101101110    1001110101101111    1001110101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40300 - 40304

  --1001110101110001    1001110101110010    1001110101110011    1001110101110100    1001110101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40305 - 40309

  --1001110101110110    1001110101110111    1001110101111000    1001110101111001    1001110101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40310 - 40314

  --1001110101111011    1001110101111100    1001110101111101    1001110101111110    1001110101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40315 - 40319

  --1001110110000000    1001110110000001    1001110110000010    1001110110000011    1001110110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40320 - 40324

  --1001110110000101    1001110110000110    1001110110000111    1001110110001000    1001110110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40325 - 40329

  --1001110110001010    1001110110001011    1001110110001100    1001110110001101    1001110110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40330 - 40334

  --1001110110001111    1001110110010000    1001110110010001    1001110110010010    1001110110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40335 - 40339

  --1001110110010100    1001110110010101    1001110110010110    1001110110010111    1001110110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40340 - 40344

  --1001110110011001    1001110110011010    1001110110011011    1001110110011100    1001110110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40345 - 40349

  --1001110110011110    1001110110011111    1001110110100000    1001110110100001    1001110110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40350 - 40354

  --1001110110100011    1001110110100100    1001110110100101    1001110110100110    1001110110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40355 - 40359

  --1001110110101000    1001110110101001    1001110110101010    1001110110101011    1001110110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40360 - 40364

  --1001110110101101    1001110110101110    1001110110101111    1001110110110000    1001110110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40365 - 40369

  --1001110110110010    1001110110110011    1001110110110100    1001110110110101    1001110110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40370 - 40374

  --1001110110110111    1001110110111000    1001110110111001    1001110110111010    1001110110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40375 - 40379

  --1001110110111100    1001110110111101    1001110110111110    1001110110111111    1001110111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40380 - 40384

  --1001110111000001    1001110111000010    1001110111000011    1001110111000100    1001110111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40385 - 40389

  --1001110111000110    1001110111000111    1001110111001000    1001110111001001    1001110111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40390 - 40394

  --1001110111001011    1001110111001100    1001110111001101    1001110111001110    1001110111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40395 - 40399

  --1001110111010000    1001110111010001    1001110111010010    1001110111010011    1001110111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40400 - 40404

  --1001110111010101    1001110111010110    1001110111010111    1001110111011000    1001110111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40405 - 40409

  --1001110111011010    1001110111011011    1001110111011100    1001110111011101    1001110111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40410 - 40414

  --1001110111011111    1001110111100000    1001110111100001    1001110111100010    1001110111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40415 - 40419

  --1001110111100100    1001110111100101    1001110111100110    1001110111100111    1001110111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40420 - 40424

  --1001110111101001    1001110111101010    1001110111101011    1001110111101100    1001110111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40425 - 40429

  --1001110111101110    1001110111101111    1001110111110000    1001110111110001    1001110111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40430 - 40434

  --1001110111110011    1001110111110100    1001110111110101    1001110111110110    1001110111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40435 - 40439

  --1001110111111000    1001110111111001    1001110111111010    1001110111111011    1001110111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40440 - 40444

  --1001110111111101    1001110111111110    1001110111111111    1001111000000000    1001111000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40445 - 40449

  --1001111000000010    1001111000000011    1001111000000100    1001111000000101    1001111000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40450 - 40454

  --1001111000000111    1001111000001000    1001111000001001    1001111000001010    1001111000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40455 - 40459

  --1001111000001100    1001111000001101    1001111000001110    1001111000001111    1001111000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40460 - 40464

  --1001111000010001    1001111000010010    1001111000010011    1001111000010100    1001111000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40465 - 40469

  --1001111000010110    1001111000010111    1001111000011000    1001111000011001    1001111000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40470 - 40474

  --1001111000011011    1001111000011100    1001111000011101    1001111000011110    1001111000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40475 - 40479

  --1001111000100000    1001111000100001    1001111000100010    1001111000100011    1001111000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40480 - 40484

  --1001111000100101    1001111000100110    1001111000100111    1001111000101000    1001111000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40485 - 40489

  --1001111000101010    1001111000101011    1001111000101100    1001111000101101    1001111000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40490 - 40494

  --1001111000101111    1001111000110000    1001111000110001    1001111000110010    1001111000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40495 - 40499

  --1001111000110100    1001111000110101    1001111000110110    1001111000110111    1001111000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40500 - 40504

  --1001111000111001    1001111000111010    1001111000111011    1001111000111100    1001111000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40505 - 40509

  --1001111000111110    1001111000111111    1001111001000000    1001111001000001    1001111001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40510 - 40514

  --1001111001000011    1001111001000100    1001111001000101    1001111001000110    1001111001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40515 - 40519

  --1001111001001000    1001111001001001    1001111001001010    1001111001001011    1001111001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40520 - 40524

  --1001111001001101    1001111001001110    1001111001001111    1001111001010000    1001111001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40525 - 40529

  --1001111001010010    1001111001010011    1001111001010100    1001111001010101    1001111001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40530 - 40534

  --1001111001010111    1001111001011000    1001111001011001    1001111001011010    1001111001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40535 - 40539

  --1001111001011100    1001111001011101    1001111001011110    1001111001011111    1001111001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40540 - 40544

  --1001111001100001    1001111001100010    1001111001100011    1001111001100100    1001111001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40545 - 40549

  --1001111001100110    1001111001100111    1001111001101000    1001111001101001    1001111001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40550 - 40554

  --1001111001101011    1001111001101100    1001111001101101    1001111001101110    1001111001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40555 - 40559

  --1001111001110000    1001111001110001    1001111001110010    1001111001110011    1001111001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40560 - 40564

  --1001111001110101    1001111001110110    1001111001110111    1001111001111000    1001111001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40565 - 40569

  --1001111001111010    1001111001111011    1001111001111100    1001111001111101    1001111001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40570 - 40574

  --1001111001111111    1001111010000000    1001111010000001    1001111010000010    1001111010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40575 - 40579

  --1001111010000100    1001111010000101    1001111010000110    1001111010000111    1001111010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40580 - 40584

  --1001111010001001    1001111010001010    1001111010001011    1001111010001100    1001111010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40585 - 40589

  --1001111010001110    1001111010001111    1001111010010000    1001111010010001    1001111010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40590 - 40594

  --1001111010010011    1001111010010100    1001111010010101    1001111010010110    1001111010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40595 - 40599

  --1001111010011000    1001111010011001    1001111010011010    1001111010011011    1001111010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40600 - 40604

  --1001111010011101    1001111010011110    1001111010011111    1001111010100000    1001111010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40605 - 40609

  --1001111010100010    1001111010100011    1001111010100100    1001111010100101    1001111010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40610 - 40614

  --1001111010100111    1001111010101000    1001111010101001    1001111010101010    1001111010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40615 - 40619

  --1001111010101100    1001111010101101    1001111010101110    1001111010101111    1001111010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40620 - 40624

  --1001111010110001    1001111010110010    1001111010110011    1001111010110100    1001111010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40625 - 40629

  --1001111010110110    1001111010110111    1001111010111000    1001111010111001    1001111010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40630 - 40634

  --1001111010111011    1001111010111100    1001111010111101    1001111010111110    1001111010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40635 - 40639

  --1001111011000000    1001111011000001    1001111011000010    1001111011000011    1001111011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40640 - 40644

  --1001111011000101    1001111011000110    1001111011000111    1001111011001000    1001111011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40645 - 40649

  --1001111011001010    1001111011001011    1001111011001100    1001111011001101    1001111011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40650 - 40654

  --1001111011001111    1001111011010000    1001111011010001    1001111011010010    1001111011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40655 - 40659

  --1001111011010100    1001111011010101    1001111011010110    1001111011010111    1001111011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40660 - 40664

  --1001111011011001    1001111011011010    1001111011011011    1001111011011100    1001111011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40665 - 40669

  --1001111011011110    1001111011011111    1001111011100000    1001111011100001    1001111011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40670 - 40674

  --1001111011100011    1001111011100100    1001111011100101    1001111011100110    1001111011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40675 - 40679

  --1001111011101000    1001111011101001    1001111011101010    1001111011101011    1001111011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40680 - 40684

  --1001111011101101    1001111011101110    1001111011101111    1001111011110000    1001111011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40685 - 40689

  --1001111011110010    1001111011110011    1001111011110100    1001111011110101    1001111011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40690 - 40694

  --1001111011110111    1001111011111000    1001111011111001    1001111011111010    1001111011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40695 - 40699

  --1001111011111100    1001111011111101    1001111011111110    1001111011111111    1001111100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40700 - 40704

  --1001111100000001    1001111100000010    1001111100000011    1001111100000100    1001111100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40705 - 40709

  --1001111100000110    1001111100000111    1001111100001000    1001111100001001    1001111100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40710 - 40714

  --1001111100001011    1001111100001100    1001111100001101    1001111100001110    1001111100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40715 - 40719

  --1001111100010000    1001111100010001    1001111100010010    1001111100010011    1001111100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40720 - 40724

  --1001111100010101    1001111100010110    1001111100010111    1001111100011000    1001111100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40725 - 40729

  --1001111100011010    1001111100011011    1001111100011100    1001111100011101    1001111100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40730 - 40734

  --1001111100011111    1001111100100000    1001111100100001    1001111100100010    1001111100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40735 - 40739

  --1001111100100100    1001111100100101    1001111100100110    1001111100100111    1001111100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40740 - 40744

  --1001111100101001    1001111100101010    1001111100101011    1001111100101100    1001111100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40745 - 40749

  --1001111100101110    1001111100101111    1001111100110000    1001111100110001    1001111100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40750 - 40754

  --1001111100110011    1001111100110100    1001111100110101    1001111100110110    1001111100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40755 - 40759

  --1001111100111000    1001111100111001    1001111100111010    1001111100111011    1001111100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40760 - 40764

  --1001111100111101    1001111100111110    1001111100111111    1001111101000000    1001111101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40765 - 40769

  --1001111101000010    1001111101000011    1001111101000100    1001111101000101    1001111101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40770 - 40774

  --1001111101000111    1001111101001000    1001111101001001    1001111101001010    1001111101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40775 - 40779

  --1001111101001100    1001111101001101    1001111101001110    1001111101001111    1001111101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40780 - 40784

  --1001111101010001    1001111101010010    1001111101010011    1001111101010100    1001111101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40785 - 40789

  --1001111101010110    1001111101010111    1001111101011000    1001111101011001    1001111101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40790 - 40794

  --1001111101011011    1001111101011100    1001111101011101    1001111101011110    1001111101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40795 - 40799

  --1001111101100000    1001111101100001    1001111101100010    1001111101100011    1001111101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40800 - 40804

  --1001111101100101    1001111101100110    1001111101100111    1001111101101000    1001111101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40805 - 40809

  --1001111101101010    1001111101101011    1001111101101100    1001111101101101    1001111101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40810 - 40814

  --1001111101101111    1001111101110000    1001111101110001    1001111101110010    1001111101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40815 - 40819

  --1001111101110100    1001111101110101    1001111101110110    1001111101110111    1001111101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40820 - 40824

  --1001111101111001    1001111101111010    1001111101111011    1001111101111100    1001111101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40825 - 40829

  --1001111101111110    1001111101111111    1001111110000000    1001111110000001    1001111110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40830 - 40834

  --1001111110000011    1001111110000100    1001111110000101    1001111110000110    1001111110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40835 - 40839

  --1001111110001000    1001111110001001    1001111110001010    1001111110001011    1001111110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40840 - 40844

  --1001111110001101    1001111110001110    1001111110001111    1001111110010000    1001111110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40845 - 40849

  --1001111110010010    1001111110010011    1001111110010100    1001111110010101    1001111110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40850 - 40854

  --1001111110010111    1001111110011000    1001111110011001    1001111110011010    1001111110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40855 - 40859

  --1001111110011100    1001111110011101    1001111110011110    1001111110011111    1001111110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40860 - 40864

  --1001111110100001    1001111110100010    1001111110100011    1001111110100100    1001111110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40865 - 40869

  --1001111110100110    1001111110100111    1001111110101000    1001111110101001    1001111110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40870 - 40874

  --1001111110101011    1001111110101100    1001111110101101    1001111110101110    1001111110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40875 - 40879

  --1001111110110000    1001111110110001    1001111110110010    1001111110110011    1001111110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40880 - 40884

  --1001111110110101    1001111110110110    1001111110110111    1001111110111000    1001111110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40885 - 40889

  --1001111110111010    1001111110111011    1001111110111100    1001111110111101    1001111110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40890 - 40894

  --1001111110111111    1001111111000000    1001111111000001    1001111111000010    1001111111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40895 - 40899

  --1001111111000100    1001111111000101    1001111111000110    1001111111000111    1001111111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40900 - 40904

  --1001111111001001    1001111111001010    1001111111001011    1001111111001100    1001111111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40905 - 40909

  --1001111111001110    1001111111001111    1001111111010000    1001111111010001    1001111111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40910 - 40914

  --1001111111010011    1001111111010100    1001111111010101    1001111111010110    1001111111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40915 - 40919

  --1001111111011000    1001111111011001    1001111111011010    1001111111011011    1001111111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40920 - 40924

  --1001111111011101    1001111111011110    1001111111011111    1001111111100000    1001111111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40925 - 40929

  --1001111111100010    1001111111100011    1001111111100100    1001111111100101    1001111111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40930 - 40934

  --1001111111100111    1001111111101000    1001111111101001    1001111111101010    1001111111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40935 - 40939

  --1001111111101100    1001111111101101    1001111111101110    1001111111101111    1001111111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40940 - 40944

  --1001111111110001    1001111111110010    1001111111110011    1001111111110100    1001111111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40945 - 40949

  --1001111111110110    1001111111110111    1001111111111000    1001111111111001    1001111111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40950 - 40954

  --1001111111111011    1001111111111100    1001111111111101    1001111111111110    1001111111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40955 - 40959

  --1010000000000000    1010000000000001    1010000000000010    1010000000000011    1010000000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40960 - 40964

  --1010000000000101    1010000000000110    1010000000000111    1010000000001000    1010000000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40965 - 40969

  --1010000000001010    1010000000001011    1010000000001100    1010000000001101    1010000000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40970 - 40974

  --1010000000001111    1010000000010000    1010000000010001    1010000000010010    1010000000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40975 - 40979

  --1010000000010100    1010000000010101    1010000000010110    1010000000010111    1010000000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40980 - 40984

  --1010000000011001    1010000000011010    1010000000011011    1010000000011100    1010000000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40985 - 40989

  --1010000000011110    1010000000011111    1010000000100000    1010000000100001    1010000000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40990 - 40994

  --1010000000100011    1010000000100100    1010000000100101    1010000000100110    1010000000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 40995 - 40999

  --1010000000101000    1010000000101001    1010000000101010    1010000000101011    1010000000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41000 - 41004

  --1010000000101101    1010000000101110    1010000000101111    1010000000110000    1010000000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41005 - 41009

  --1010000000110010    1010000000110011    1010000000110100    1010000000110101    1010000000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41010 - 41014

  --1010000000110111    1010000000111000    1010000000111001    1010000000111010    1010000000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41015 - 41019

  --1010000000111100    1010000000111101    1010000000111110    1010000000111111    1010000001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41020 - 41024

  --1010000001000001    1010000001000010    1010000001000011    1010000001000100    1010000001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41025 - 41029

  --1010000001000110    1010000001000111    1010000001001000    1010000001001001    1010000001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41030 - 41034

  --1010000001001011    1010000001001100    1010000001001101    1010000001001110    1010000001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41035 - 41039

  --1010000001010000    1010000001010001    1010000001010010    1010000001010011    1010000001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41040 - 41044

  --1010000001010101    1010000001010110    1010000001010111    1010000001011000    1010000001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41045 - 41049

  --1010000001011010    1010000001011011    1010000001011100    1010000001011101    1010000001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41050 - 41054

  --1010000001011111    1010000001100000    1010000001100001    1010000001100010    1010000001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41055 - 41059

  --1010000001100100    1010000001100101    1010000001100110    1010000001100111    1010000001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41060 - 41064

  --1010000001101001    1010000001101010    1010000001101011    1010000001101100    1010000001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41065 - 41069

  --1010000001101110    1010000001101111    1010000001110000    1010000001110001    1010000001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41070 - 41074

  --1010000001110011    1010000001110100    1010000001110101    1010000001110110    1010000001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41075 - 41079

  --1010000001111000    1010000001111001    1010000001111010    1010000001111011    1010000001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41080 - 41084

  --1010000001111101    1010000001111110    1010000001111111    1010000010000000    1010000010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41085 - 41089

  --1010000010000010    1010000010000011    1010000010000100    1010000010000101    1010000010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41090 - 41094

  --1010000010000111    1010000010001000    1010000010001001    1010000010001010    1010000010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41095 - 41099

  --1010000010001100    1010000010001101    1010000010001110    1010000010001111    1010000010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41100 - 41104

  --1010000010010001    1010000010010010    1010000010010011    1010000010010100    1010000010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41105 - 41109

  --1010000010010110    1010000010010111    1010000010011000    1010000010011001    1010000010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41110 - 41114

  --1010000010011011    1010000010011100    1010000010011101    1010000010011110    1010000010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41115 - 41119

  --1010000010100000    1010000010100001    1010000010100010    1010000010100011    1010000010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41120 - 41124

  --1010000010100101    1010000010100110    1010000010100111    1010000010101000    1010000010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41125 - 41129

  --1010000010101010    1010000010101011    1010000010101100    1010000010101101    1010000010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41130 - 41134

  --1010000010101111    1010000010110000    1010000010110001    1010000010110010    1010000010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41135 - 41139

  --1010000010110100    1010000010110101    1010000010110110    1010000010110111    1010000010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41140 - 41144

  --1010000010111001    1010000010111010    1010000010111011    1010000010111100    1010000010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41145 - 41149

  --1010000010111110    1010000010111111    1010000011000000    1010000011000001    1010000011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41150 - 41154

  --1010000011000011    1010000011000100    1010000011000101    1010000011000110    1010000011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41155 - 41159

  --1010000011001000    1010000011001001    1010000011001010    1010000011001011    1010000011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41160 - 41164

  --1010000011001101    1010000011001110    1010000011001111    1010000011010000    1010000011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41165 - 41169

  --1010000011010010    1010000011010011    1010000011010100    1010000011010101    1010000011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41170 - 41174

  --1010000011010111    1010000011011000    1010000011011001    1010000011011010    1010000011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41175 - 41179

  --1010000011011100    1010000011011101    1010000011011110    1010000011011111    1010000011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41180 - 41184

  --1010000011100001    1010000011100010    1010000011100011    1010000011100100    1010000011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41185 - 41189

  --1010000011100110    1010000011100111    1010000011101000    1010000011101001    1010000011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41190 - 41194

  --1010000011101011    1010000011101100    1010000011101101    1010000011101110    1010000011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41195 - 41199

  --1010000011110000    1010000011110001    1010000011110010    1010000011110011    1010000011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41200 - 41204

  --1010000011110101    1010000011110110    1010000011110111    1010000011111000    1010000011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41205 - 41209

  --1010000011111010    1010000011111011    1010000011111100    1010000011111101    1010000011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41210 - 41214

  --1010000011111111    1010000100000000    1010000100000001    1010000100000010    1010000100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41215 - 41219

  --1010000100000100    1010000100000101    1010000100000110    1010000100000111    1010000100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41220 - 41224

  --1010000100001001    1010000100001010    1010000100001011    1010000100001100    1010000100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41225 - 41229

  --1010000100001110    1010000100001111    1010000100010000    1010000100010001    1010000100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41230 - 41234

  --1010000100010011    1010000100010100    1010000100010101    1010000100010110    1010000100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41235 - 41239

  --1010000100011000    1010000100011001    1010000100011010    1010000100011011    1010000100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41240 - 41244

  --1010000100011101    1010000100011110    1010000100011111    1010000100100000    1010000100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41245 - 41249

  --1010000100100010    1010000100100011    1010000100100100    1010000100100101    1010000100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41250 - 41254

  --1010000100100111    1010000100101000    1010000100101001    1010000100101010    1010000100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41255 - 41259

  --1010000100101100    1010000100101101    1010000100101110    1010000100101111    1010000100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41260 - 41264

  --1010000100110001    1010000100110010    1010000100110011    1010000100110100    1010000100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41265 - 41269

  --1010000100110110    1010000100110111    1010000100111000    1010000100111001    1010000100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41270 - 41274

  --1010000100111011    1010000100111100    1010000100111101    1010000100111110    1010000100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41275 - 41279

  --1010000101000000    1010000101000001    1010000101000010    1010000101000011    1010000101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41280 - 41284

  --1010000101000101    1010000101000110    1010000101000111    1010000101001000    1010000101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41285 - 41289

  --1010000101001010    1010000101001011    1010000101001100    1010000101001101    1010000101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41290 - 41294

  --1010000101001111    1010000101010000    1010000101010001    1010000101010010    1010000101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41295 - 41299

  --1010000101010100    1010000101010101    1010000101010110    1010000101010111    1010000101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41300 - 41304

  --1010000101011001    1010000101011010    1010000101011011    1010000101011100    1010000101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41305 - 41309

  --1010000101011110    1010000101011111    1010000101100000    1010000101100001    1010000101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41310 - 41314

  --1010000101100011    1010000101100100    1010000101100101    1010000101100110    1010000101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41315 - 41319

  --1010000101101000    1010000101101001    1010000101101010    1010000101101011    1010000101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41320 - 41324

  --1010000101101101    1010000101101110    1010000101101111    1010000101110000    1010000101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41325 - 41329

  --1010000101110010    1010000101110011    1010000101110100    1010000101110101    1010000101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41330 - 41334

  --1010000101110111    1010000101111000    1010000101111001    1010000101111010    1010000101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41335 - 41339

  --1010000101111100    1010000101111101    1010000101111110    1010000101111111    1010000110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41340 - 41344

  --1010000110000001    1010000110000010    1010000110000011    1010000110000100    1010000110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41345 - 41349

  --1010000110000110    1010000110000111    1010000110001000    1010000110001001    1010000110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41350 - 41354

  --1010000110001011    1010000110001100    1010000110001101    1010000110001110    1010000110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41355 - 41359

  --1010000110010000    1010000110010001    1010000110010010    1010000110010011    1010000110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41360 - 41364

  --1010000110010101    1010000110010110    1010000110010111    1010000110011000    1010000110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41365 - 41369

  --1010000110011010    1010000110011011    1010000110011100    1010000110011101    1010000110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41370 - 41374

  --1010000110011111    1010000110100000    1010000110100001    1010000110100010    1010000110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41375 - 41379

  --1010000110100100    1010000110100101    1010000110100110    1010000110100111    1010000110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41380 - 41384

  --1010000110101001    1010000110101010    1010000110101011    1010000110101100    1010000110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41385 - 41389

  --1010000110101110    1010000110101111    1010000110110000    1010000110110001    1010000110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41390 - 41394

  --1010000110110011    1010000110110100    1010000110110101    1010000110110110    1010000110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41395 - 41399

  --1010000110111000    1010000110111001    1010000110111010    1010000110111011    1010000110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41400 - 41404

  --1010000110111101    1010000110111110    1010000110111111    1010000111000000    1010000111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41405 - 41409

  --1010000111000010    1010000111000011    1010000111000100    1010000111000101    1010000111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41410 - 41414

  --1010000111000111    1010000111001000    1010000111001001    1010000111001010    1010000111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41415 - 41419

  --1010000111001100    1010000111001101    1010000111001110    1010000111001111    1010000111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41420 - 41424

  --1010000111010001    1010000111010010    1010000111010011    1010000111010100    1010000111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41425 - 41429

  --1010000111010110    1010000111010111    1010000111011000    1010000111011001    1010000111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41430 - 41434

  --1010000111011011    1010000111011100    1010000111011101    1010000111011110    1010000111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41435 - 41439

  --1010000111100000    1010000111100001    1010000111100010    1010000111100011    1010000111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41440 - 41444

  --1010000111100101    1010000111100110    1010000111100111    1010000111101000    1010000111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41445 - 41449

  --1010000111101010    1010000111101011    1010000111101100    1010000111101101    1010000111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41450 - 41454

  --1010000111101111    1010000111110000    1010000111110001    1010000111110010    1010000111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41455 - 41459

  --1010000111110100    1010000111110101    1010000111110110    1010000111110111    1010000111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41460 - 41464

  --1010000111111001    1010000111111010    1010000111111011    1010000111111100    1010000111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41465 - 41469

  --1010000111111110    1010000111111111    1010001000000000    1010001000000001    1010001000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41470 - 41474

  --1010001000000011    1010001000000100    1010001000000101    1010001000000110    1010001000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41475 - 41479

  --1010001000001000    1010001000001001    1010001000001010    1010001000001011    1010001000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41480 - 41484

  --1010001000001101    1010001000001110    1010001000001111    1010001000010000    1010001000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41485 - 41489

  --1010001000010010    1010001000010011    1010001000010100    1010001000010101    1010001000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41490 - 41494

  --1010001000010111    1010001000011000    1010001000011001    1010001000011010    1010001000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41495 - 41499

  --1010001000011100    1010001000011101    1010001000011110    1010001000011111    1010001000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41500 - 41504

  --1010001000100001    1010001000100010    1010001000100011    1010001000100100    1010001000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41505 - 41509

  --1010001000100110    1010001000100111    1010001000101000    1010001000101001    1010001000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41510 - 41514

  --1010001000101011    1010001000101100    1010001000101101    1010001000101110    1010001000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41515 - 41519

  --1010001000110000    1010001000110001    1010001000110010    1010001000110011    1010001000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41520 - 41524

  --1010001000110101    1010001000110110    1010001000110111    1010001000111000    1010001000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41525 - 41529

  --1010001000111010    1010001000111011    1010001000111100    1010001000111101    1010001000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41530 - 41534

  --1010001000111111    1010001001000000    1010001001000001    1010001001000010    1010001001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41535 - 41539

  --1010001001000100    1010001001000101    1010001001000110    1010001001000111    1010001001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41540 - 41544

  --1010001001001001    1010001001001010    1010001001001011    1010001001001100    1010001001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41545 - 41549

  --1010001001001110    1010001001001111    1010001001010000    1010001001010001    1010001001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41550 - 41554

  --1010001001010011    1010001001010100    1010001001010101    1010001001010110    1010001001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41555 - 41559

  --1010001001011000    1010001001011001    1010001001011010    1010001001011011    1010001001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41560 - 41564

  --1010001001011101    1010001001011110    1010001001011111    1010001001100000    1010001001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41565 - 41569

  --1010001001100010    1010001001100011    1010001001100100    1010001001100101    1010001001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41570 - 41574

  --1010001001100111    1010001001101000    1010001001101001    1010001001101010    1010001001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41575 - 41579

  --1010001001101100    1010001001101101    1010001001101110    1010001001101111    1010001001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41580 - 41584

  --1010001001110001    1010001001110010    1010001001110011    1010001001110100    1010001001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41585 - 41589

  --1010001001110110    1010001001110111    1010001001111000    1010001001111001    1010001001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41590 - 41594

  --1010001001111011    1010001001111100    1010001001111101    1010001001111110    1010001001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41595 - 41599

  --1010001010000000    1010001010000001    1010001010000010    1010001010000011    1010001010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41600 - 41604

  --1010001010000101    1010001010000110    1010001010000111    1010001010001000    1010001010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41605 - 41609

  --1010001010001010    1010001010001011    1010001010001100    1010001010001101    1010001010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41610 - 41614

  --1010001010001111    1010001010010000    1010001010010001    1010001010010010    1010001010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41615 - 41619

  --1010001010010100    1010001010010101    1010001010010110    1010001010010111    1010001010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41620 - 41624

  --1010001010011001    1010001010011010    1010001010011011    1010001010011100    1010001010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41625 - 41629

  --1010001010011110    1010001010011111    1010001010100000    1010001010100001    1010001010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41630 - 41634

  --1010001010100011    1010001010100100    1010001010100101    1010001010100110    1010001010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41635 - 41639

  --1010001010101000    1010001010101001    1010001010101010    1010001010101011    1010001010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41640 - 41644

  --1010001010101101    1010001010101110    1010001010101111    1010001010110000    1010001010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41645 - 41649

  --1010001010110010    1010001010110011    1010001010110100    1010001010110101    1010001010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41650 - 41654

  --1010001010110111    1010001010111000    1010001010111001    1010001010111010    1010001010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41655 - 41659

  --1010001010111100    1010001010111101    1010001010111110    1010001010111111    1010001011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41660 - 41664

  --1010001011000001    1010001011000010    1010001011000011    1010001011000100    1010001011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41665 - 41669

  --1010001011000110    1010001011000111    1010001011001000    1010001011001001    1010001011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41670 - 41674

  --1010001011001011    1010001011001100    1010001011001101    1010001011001110    1010001011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41675 - 41679

  --1010001011010000    1010001011010001    1010001011010010    1010001011010011    1010001011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41680 - 41684

  --1010001011010101    1010001011010110    1010001011010111    1010001011011000    1010001011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41685 - 41689

  --1010001011011010    1010001011011011    1010001011011100    1010001011011101    1010001011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41690 - 41694

  --1010001011011111    1010001011100000    1010001011100001    1010001011100010    1010001011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41695 - 41699

  --1010001011100100    1010001011100101    1010001011100110    1010001011100111    1010001011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41700 - 41704

  --1010001011101001    1010001011101010    1010001011101011    1010001011101100    1010001011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41705 - 41709

  --1010001011101110    1010001011101111    1010001011110000    1010001011110001    1010001011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41710 - 41714

  --1010001011110011    1010001011110100    1010001011110101    1010001011110110    1010001011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41715 - 41719

  --1010001011111000    1010001011111001    1010001011111010    1010001011111011    1010001011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41720 - 41724

  --1010001011111101    1010001011111110    1010001011111111    1010001100000000    1010001100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41725 - 41729

  --1010001100000010    1010001100000011    1010001100000100    1010001100000101    1010001100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41730 - 41734

  --1010001100000111    1010001100001000    1010001100001001    1010001100001010    1010001100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41735 - 41739

  --1010001100001100    1010001100001101    1010001100001110    1010001100001111    1010001100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41740 - 41744

  --1010001100010001    1010001100010010    1010001100010011    1010001100010100    1010001100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41745 - 41749

  --1010001100010110    1010001100010111    1010001100011000    1010001100011001    1010001100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41750 - 41754

  --1010001100011011    1010001100011100    1010001100011101    1010001100011110    1010001100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41755 - 41759

  --1010001100100000    1010001100100001    1010001100100010    1010001100100011    1010001100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41760 - 41764

  --1010001100100101    1010001100100110    1010001100100111    1010001100101000    1010001100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41765 - 41769

  --1010001100101010    1010001100101011    1010001100101100    1010001100101101    1010001100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41770 - 41774

  --1010001100101111    1010001100110000    1010001100110001    1010001100110010    1010001100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41775 - 41779

  --1010001100110100    1010001100110101    1010001100110110    1010001100110111    1010001100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41780 - 41784

  --1010001100111001    1010001100111010    1010001100111011    1010001100111100    1010001100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41785 - 41789

  --1010001100111110    1010001100111111    1010001101000000    1010001101000001    1010001101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41790 - 41794

  --1010001101000011    1010001101000100    1010001101000101    1010001101000110    1010001101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41795 - 41799

  --1010001101001000    1010001101001001    1010001101001010    1010001101001011    1010001101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41800 - 41804

  --1010001101001101    1010001101001110    1010001101001111    1010001101010000    1010001101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41805 - 41809

  --1010001101010010    1010001101010011    1010001101010100    1010001101010101    1010001101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41810 - 41814

  --1010001101010111    1010001101011000    1010001101011001    1010001101011010    1010001101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41815 - 41819

  --1010001101011100    1010001101011101    1010001101011110    1010001101011111    1010001101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41820 - 41824

  --1010001101100001    1010001101100010    1010001101100011    1010001101100100    1010001101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41825 - 41829

  --1010001101100110    1010001101100111    1010001101101000    1010001101101001    1010001101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41830 - 41834

  --1010001101101011    1010001101101100    1010001101101101    1010001101101110    1010001101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41835 - 41839

  --1010001101110000    1010001101110001    1010001101110010    1010001101110011    1010001101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41840 - 41844

  --1010001101110101    1010001101110110    1010001101110111    1010001101111000    1010001101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41845 - 41849

  --1010001101111010    1010001101111011    1010001101111100    1010001101111101    1010001101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41850 - 41854

  --1010001101111111    1010001110000000    1010001110000001    1010001110000010    1010001110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41855 - 41859

  --1010001110000100    1010001110000101    1010001110000110    1010001110000111    1010001110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41860 - 41864

  --1010001110001001    1010001110001010    1010001110001011    1010001110001100    1010001110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41865 - 41869

  --1010001110001110    1010001110001111    1010001110010000    1010001110010001    1010001110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41870 - 41874

  --1010001110010011    1010001110010100    1010001110010101    1010001110010110    1010001110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41875 - 41879

  --1010001110011000    1010001110011001    1010001110011010    1010001110011011    1010001110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41880 - 41884

  --1010001110011101    1010001110011110    1010001110011111    1010001110100000    1010001110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41885 - 41889

  --1010001110100010    1010001110100011    1010001110100100    1010001110100101    1010001110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41890 - 41894

  --1010001110100111    1010001110101000    1010001110101001    1010001110101010    1010001110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41895 - 41899

  --1010001110101100    1010001110101101    1010001110101110    1010001110101111    1010001110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41900 - 41904

  --1010001110110001    1010001110110010    1010001110110011    1010001110110100    1010001110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41905 - 41909

  --1010001110110110    1010001110110111    1010001110111000    1010001110111001    1010001110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41910 - 41914

  --1010001110111011    1010001110111100    1010001110111101    1010001110111110    1010001110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41915 - 41919

  --1010001111000000    1010001111000001    1010001111000010    1010001111000011    1010001111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41920 - 41924

  --1010001111000101    1010001111000110    1010001111000111    1010001111001000    1010001111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41925 - 41929

  --1010001111001010    1010001111001011    1010001111001100    1010001111001101    1010001111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41930 - 41934

  --1010001111001111    1010001111010000    1010001111010001    1010001111010010    1010001111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41935 - 41939

  --1010001111010100    1010001111010101    1010001111010110    1010001111010111    1010001111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41940 - 41944

  --1010001111011001    1010001111011010    1010001111011011    1010001111011100    1010001111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41945 - 41949

  --1010001111011110    1010001111011111    1010001111100000    1010001111100001    1010001111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41950 - 41954

  --1010001111100011    1010001111100100    1010001111100101    1010001111100110    1010001111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41955 - 41959

  --1010001111101000    1010001111101001    1010001111101010    1010001111101011    1010001111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41960 - 41964

  --1010001111101101    1010001111101110    1010001111101111    1010001111110000    1010001111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41965 - 41969

  --1010001111110010    1010001111110011    1010001111110100    1010001111110101    1010001111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41970 - 41974

  --1010001111110111    1010001111111000    1010001111111001    1010001111111010    1010001111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41975 - 41979

  --1010001111111100    1010001111111101    1010001111111110    1010001111111111    1010010000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41980 - 41984

  --1010010000000001    1010010000000010    1010010000000011    1010010000000100    1010010000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41985 - 41989

  --1010010000000110    1010010000000111    1010010000001000    1010010000001001    1010010000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41990 - 41994

  --1010010000001011    1010010000001100    1010010000001101    1010010000001110    1010010000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 41995 - 41999

  --1010010000010000    1010010000010001    1010010000010010    1010010000010011    1010010000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42000 - 42004

  --1010010000010101    1010010000010110    1010010000010111    1010010000011000    1010010000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42005 - 42009

  --1010010000011010    1010010000011011    1010010000011100    1010010000011101    1010010000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42010 - 42014

  --1010010000011111    1010010000100000    1010010000100001    1010010000100010    1010010000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42015 - 42019

  --1010010000100100    1010010000100101    1010010000100110    1010010000100111    1010010000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42020 - 42024

  --1010010000101001    1010010000101010    1010010000101011    1010010000101100    1010010000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42025 - 42029

  --1010010000101110    1010010000101111    1010010000110000    1010010000110001    1010010000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42030 - 42034

  --1010010000110011    1010010000110100    1010010000110101    1010010000110110    1010010000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42035 - 42039

  --1010010000111000    1010010000111001    1010010000111010    1010010000111011    1010010000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42040 - 42044

  --1010010000111101    1010010000111110    1010010000111111    1010010001000000    1010010001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42045 - 42049

  --1010010001000010    1010010001000011    1010010001000100    1010010001000101    1010010001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42050 - 42054

  --1010010001000111    1010010001001000    1010010001001001    1010010001001010    1010010001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42055 - 42059

  --1010010001001100    1010010001001101    1010010001001110    1010010001001111    1010010001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42060 - 42064

  --1010010001010001    1010010001010010    1010010001010011    1010010001010100    1010010001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42065 - 42069

  --1010010001010110    1010010001010111    1010010001011000    1010010001011001    1010010001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42070 - 42074

  --1010010001011011    1010010001011100    1010010001011101    1010010001011110    1010010001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42075 - 42079

  --1010010001100000    1010010001100001    1010010001100010    1010010001100011    1010010001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42080 - 42084

  --1010010001100101    1010010001100110    1010010001100111    1010010001101000    1010010001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42085 - 42089

  --1010010001101010    1010010001101011    1010010001101100    1010010001101101    1010010001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42090 - 42094

  --1010010001101111    1010010001110000    1010010001110001    1010010001110010    1010010001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42095 - 42099

  --1010010001110100    1010010001110101    1010010001110110    1010010001110111    1010010001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42100 - 42104

  --1010010001111001    1010010001111010    1010010001111011    1010010001111100    1010010001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42105 - 42109

  --1010010001111110    1010010001111111    1010010010000000    1010010010000001    1010010010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42110 - 42114

  --1010010010000011    1010010010000100    1010010010000101    1010010010000110    1010010010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42115 - 42119

  --1010010010001000    1010010010001001    1010010010001010    1010010010001011    1010010010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42120 - 42124

  --1010010010001101    1010010010001110    1010010010001111    1010010010010000    1010010010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42125 - 42129

  --1010010010010010    1010010010010011    1010010010010100    1010010010010101    1010010010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42130 - 42134

  --1010010010010111    1010010010011000    1010010010011001    1010010010011010    1010010010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42135 - 42139

  --1010010010011100    1010010010011101    1010010010011110    1010010010011111    1010010010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42140 - 42144

  --1010010010100001    1010010010100010    1010010010100011    1010010010100100    1010010010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42145 - 42149

  --1010010010100110    1010010010100111    1010010010101000    1010010010101001    1010010010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42150 - 42154

  --1010010010101011    1010010010101100    1010010010101101    1010010010101110    1010010010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42155 - 42159

  --1010010010110000    1010010010110001    1010010010110010    1010010010110011    1010010010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42160 - 42164

  --1010010010110101    1010010010110110    1010010010110111    1010010010111000    1010010010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42165 - 42169

  --1010010010111010    1010010010111011    1010010010111100    1010010010111101    1010010010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42170 - 42174

  --1010010010111111    1010010011000000    1010010011000001    1010010011000010    1010010011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42175 - 42179

  --1010010011000100    1010010011000101    1010010011000110    1010010011000111    1010010011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42180 - 42184

  --1010010011001001    1010010011001010    1010010011001011    1010010011001100    1010010011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42185 - 42189

  --1010010011001110    1010010011001111    1010010011010000    1010010011010001    1010010011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42190 - 42194

  --1010010011010011    1010010011010100    1010010011010101    1010010011010110    1010010011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42195 - 42199

  --1010010011011000    1010010011011001    1010010011011010    1010010011011011    1010010011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42200 - 42204

  --1010010011011101    1010010011011110    1010010011011111    1010010011100000    1010010011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42205 - 42209

  --1010010011100010    1010010011100011    1010010011100100    1010010011100101    1010010011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42210 - 42214

  --1010010011100111    1010010011101000    1010010011101001    1010010011101010    1010010011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42215 - 42219

  --1010010011101100    1010010011101101    1010010011101110    1010010011101111    1010010011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42220 - 42224

  --1010010011110001    1010010011110010    1010010011110011    1010010011110100    1010010011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42225 - 42229

  --1010010011110110    1010010011110111    1010010011111000    1010010011111001    1010010011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42230 - 42234

  --1010010011111011    1010010011111100    1010010011111101    1010010011111110    1010010011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42235 - 42239

  --1010010100000000    1010010100000001    1010010100000010    1010010100000011    1010010100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42240 - 42244

  --1010010100000101    1010010100000110    1010010100000111    1010010100001000    1010010100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42245 - 42249

  --1010010100001010    1010010100001011    1010010100001100    1010010100001101    1010010100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42250 - 42254

  --1010010100001111    1010010100010000    1010010100010001    1010010100010010    1010010100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42255 - 42259

  --1010010100010100    1010010100010101    1010010100010110    1010010100010111    1010010100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42260 - 42264

  --1010010100011001    1010010100011010    1010010100011011    1010010100011100    1010010100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42265 - 42269

  --1010010100011110    1010010100011111    1010010100100000    1010010100100001    1010010100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42270 - 42274

  --1010010100100011    1010010100100100    1010010100100101    1010010100100110    1010010100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42275 - 42279

  --1010010100101000    1010010100101001    1010010100101010    1010010100101011    1010010100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42280 - 42284

  --1010010100101101    1010010100101110    1010010100101111    1010010100110000    1010010100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42285 - 42289

  --1010010100110010    1010010100110011    1010010100110100    1010010100110101    1010010100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42290 - 42294

  --1010010100110111    1010010100111000    1010010100111001    1010010100111010    1010010100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42295 - 42299

  --1010010100111100    1010010100111101    1010010100111110    1010010100111111    1010010101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42300 - 42304

  --1010010101000001    1010010101000010    1010010101000011    1010010101000100    1010010101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42305 - 42309

  --1010010101000110    1010010101000111    1010010101001000    1010010101001001    1010010101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42310 - 42314

  --1010010101001011    1010010101001100    1010010101001101    1010010101001110    1010010101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42315 - 42319

  --1010010101010000    1010010101010001    1010010101010010    1010010101010011    1010010101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42320 - 42324

  --1010010101010101    1010010101010110    1010010101010111    1010010101011000    1010010101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42325 - 42329

  --1010010101011010    1010010101011011    1010010101011100    1010010101011101    1010010101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42330 - 42334

  --1010010101011111    1010010101100000    1010010101100001    1010010101100010    1010010101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42335 - 42339

  --1010010101100100    1010010101100101    1010010101100110    1010010101100111    1010010101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42340 - 42344

  --1010010101101001    1010010101101010    1010010101101011    1010010101101100    1010010101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42345 - 42349

  --1010010101101110    1010010101101111    1010010101110000    1010010101110001    1010010101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42350 - 42354

  --1010010101110011    1010010101110100    1010010101110101    1010010101110110    1010010101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42355 - 42359

  --1010010101111000    1010010101111001    1010010101111010    1010010101111011    1010010101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42360 - 42364

  --1010010101111101    1010010101111110    1010010101111111    1010010110000000    1010010110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42365 - 42369

  --1010010110000010    1010010110000011    1010010110000100    1010010110000101    1010010110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42370 - 42374

  --1010010110000111    1010010110001000    1010010110001001    1010010110001010    1010010110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42375 - 42379

  --1010010110001100    1010010110001101    1010010110001110    1010010110001111    1010010110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42380 - 42384

  --1010010110010001    1010010110010010    1010010110010011    1010010110010100    1010010110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42385 - 42389

  --1010010110010110    1010010110010111    1010010110011000    1010010110011001    1010010110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42390 - 42394

  --1010010110011011    1010010110011100    1010010110011101    1010010110011110    1010010110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42395 - 42399

  --1010010110100000    1010010110100001    1010010110100010    1010010110100011    1010010110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42400 - 42404

  --1010010110100101    1010010110100110    1010010110100111    1010010110101000    1010010110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42405 - 42409

  --1010010110101010    1010010110101011    1010010110101100    1010010110101101    1010010110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42410 - 42414

  --1010010110101111    1010010110110000    1010010110110001    1010010110110010    1010010110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42415 - 42419

  --1010010110110100    1010010110110101    1010010110110110    1010010110110111    1010010110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42420 - 42424

  --1010010110111001    1010010110111010    1010010110111011    1010010110111100    1010010110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42425 - 42429

  --1010010110111110    1010010110111111    1010010111000000    1010010111000001    1010010111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42430 - 42434

  --1010010111000011    1010010111000100    1010010111000101    1010010111000110    1010010111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42435 - 42439

  --1010010111001000    1010010111001001    1010010111001010    1010010111001011    1010010111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42440 - 42444

  --1010010111001101    1010010111001110    1010010111001111    1010010111010000    1010010111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42445 - 42449

  --1010010111010010    1010010111010011    1010010111010100    1010010111010101    1010010111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42450 - 42454

  --1010010111010111    1010010111011000    1010010111011001    1010010111011010    1010010111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42455 - 42459

  --1010010111011100    1010010111011101    1010010111011110    1010010111011111    1010010111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42460 - 42464

  --1010010111100001    1010010111100010    1010010111100011    1010010111100100    1010010111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42465 - 42469

  --1010010111100110    1010010111100111    1010010111101000    1010010111101001    1010010111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42470 - 42474

  --1010010111101011    1010010111101100    1010010111101101    1010010111101110    1010010111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42475 - 42479

  --1010010111110000    1010010111110001    1010010111110010    1010010111110011    1010010111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42480 - 42484

  --1010010111110101    1010010111110110    1010010111110111    1010010111111000    1010010111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42485 - 42489

  --1010010111111010    1010010111111011    1010010111111100    1010010111111101    1010010111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42490 - 42494

  --1010010111111111    1010011000000000    1010011000000001    1010011000000010    1010011000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42495 - 42499

  --1010011000000100    1010011000000101    1010011000000110    1010011000000111    1010011000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42500 - 42504

  --1010011000001001    1010011000001010    1010011000001011    1010011000001100    1010011000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42505 - 42509

  --1010011000001110    1010011000001111    1010011000010000    1010011000010001    1010011000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42510 - 42514

  --1010011000010011    1010011000010100    1010011000010101    1010011000010110    1010011000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42515 - 42519

  --1010011000011000    1010011000011001    1010011000011010    1010011000011011    1010011000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42520 - 42524

  --1010011000011101    1010011000011110    1010011000011111    1010011000100000    1010011000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42525 - 42529

  --1010011000100010    1010011000100011    1010011000100100    1010011000100101    1010011000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42530 - 42534

  --1010011000100111    1010011000101000    1010011000101001    1010011000101010    1010011000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42535 - 42539

  --1010011000101100    1010011000101101    1010011000101110    1010011000101111    1010011000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42540 - 42544

  --1010011000110001    1010011000110010    1010011000110011    1010011000110100    1010011000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42545 - 42549

  --1010011000110110    1010011000110111    1010011000111000    1010011000111001    1010011000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42550 - 42554

  --1010011000111011    1010011000111100    1010011000111101    1010011000111110    1010011000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42555 - 42559

  --1010011001000000    1010011001000001    1010011001000010    1010011001000011    1010011001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42560 - 42564

  --1010011001000101    1010011001000110    1010011001000111    1010011001001000    1010011001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42565 - 42569

  --1010011001001010    1010011001001011    1010011001001100    1010011001001101    1010011001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42570 - 42574

  --1010011001001111    1010011001010000    1010011001010001    1010011001010010    1010011001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42575 - 42579

  --1010011001010100    1010011001010101    1010011001010110    1010011001010111    1010011001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42580 - 42584

  --1010011001011001    1010011001011010    1010011001011011    1010011001011100    1010011001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42585 - 42589

  --1010011001011110    1010011001011111    1010011001100000    1010011001100001    1010011001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42590 - 42594

  --1010011001100011    1010011001100100    1010011001100101    1010011001100110    1010011001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42595 - 42599

  --1010011001101000    1010011001101001    1010011001101010    1010011001101011    1010011001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42600 - 42604

  --1010011001101101    1010011001101110    1010011001101111    1010011001110000    1010011001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42605 - 42609

  --1010011001110010    1010011001110011    1010011001110100    1010011001110101    1010011001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42610 - 42614

  --1010011001110111    1010011001111000    1010011001111001    1010011001111010    1010011001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42615 - 42619

  --1010011001111100    1010011001111101    1010011001111110    1010011001111111    1010011010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42620 - 42624

  --1010011010000001    1010011010000010    1010011010000011    1010011010000100    1010011010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42625 - 42629

  --1010011010000110    1010011010000111    1010011010001000    1010011010001001    1010011010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42630 - 42634

  --1010011010001011    1010011010001100    1010011010001101    1010011010001110    1010011010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42635 - 42639

  --1010011010010000    1010011010010001    1010011010010010    1010011010010011    1010011010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42640 - 42644

  --1010011010010101    1010011010010110    1010011010010111    1010011010011000    1010011010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42645 - 42649

  --1010011010011010    1010011010011011    1010011010011100    1010011010011101    1010011010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42650 - 42654

  --1010011010011111    1010011010100000    1010011010100001    1010011010100010    1010011010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42655 - 42659

  --1010011010100100    1010011010100101    1010011010100110    1010011010100111    1010011010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42660 - 42664

  --1010011010101001    1010011010101010    1010011010101011    1010011010101100    1010011010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42665 - 42669

  --1010011010101110    1010011010101111    1010011010110000    1010011010110001    1010011010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42670 - 42674

  --1010011010110011    1010011010110100    1010011010110101    1010011010110110    1010011010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42675 - 42679

  --1010011010111000    1010011010111001    1010011010111010    1010011010111011    1010011010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42680 - 42684

  --1010011010111101    1010011010111110    1010011010111111    1010011011000000    1010011011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42685 - 42689

  --1010011011000010    1010011011000011    1010011011000100    1010011011000101    1010011011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42690 - 42694

  --1010011011000111    1010011011001000    1010011011001001    1010011011001010    1010011011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42695 - 42699

  --1010011011001100    1010011011001101    1010011011001110    1010011011001111    1010011011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42700 - 42704

  --1010011011010001    1010011011010010    1010011011010011    1010011011010100    1010011011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42705 - 42709

  --1010011011010110    1010011011010111    1010011011011000    1010011011011001    1010011011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42710 - 42714

  --1010011011011011    1010011011011100    1010011011011101    1010011011011110    1010011011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42715 - 42719

  --1010011011100000    1010011011100001    1010011011100010    1010011011100011    1010011011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42720 - 42724

  --1010011011100101    1010011011100110    1010011011100111    1010011011101000    1010011011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42725 - 42729

  --1010011011101010    1010011011101011    1010011011101100    1010011011101101    1010011011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42730 - 42734

  --1010011011101111    1010011011110000    1010011011110001    1010011011110010    1010011011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42735 - 42739

  --1010011011110100    1010011011110101    1010011011110110    1010011011110111    1010011011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42740 - 42744

  --1010011011111001    1010011011111010    1010011011111011    1010011011111100    1010011011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42745 - 42749

  --1010011011111110    1010011011111111    1010011100000000    1010011100000001    1010011100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42750 - 42754

  --1010011100000011    1010011100000100    1010011100000101    1010011100000110    1010011100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42755 - 42759

  --1010011100001000    1010011100001001    1010011100001010    1010011100001011    1010011100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42760 - 42764

  --1010011100001101    1010011100001110    1010011100001111    1010011100010000    1010011100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42765 - 42769

  --1010011100010010    1010011100010011    1010011100010100    1010011100010101    1010011100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42770 - 42774

  --1010011100010111    1010011100011000    1010011100011001    1010011100011010    1010011100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42775 - 42779

  --1010011100011100    1010011100011101    1010011100011110    1010011100011111    1010011100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42780 - 42784

  --1010011100100001    1010011100100010    1010011100100011    1010011100100100    1010011100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42785 - 42789

  --1010011100100110    1010011100100111    1010011100101000    1010011100101001    1010011100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42790 - 42794

  --1010011100101011    1010011100101100    1010011100101101    1010011100101110    1010011100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42795 - 42799

  --1010011100110000    1010011100110001    1010011100110010    1010011100110011    1010011100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42800 - 42804

  --1010011100110101    1010011100110110    1010011100110111    1010011100111000    1010011100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42805 - 42809

  --1010011100111010    1010011100111011    1010011100111100    1010011100111101    1010011100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42810 - 42814

  --1010011100111111    1010011101000000    1010011101000001    1010011101000010    1010011101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42815 - 42819

  --1010011101000100    1010011101000101    1010011101000110    1010011101000111    1010011101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42820 - 42824

  --1010011101001001    1010011101001010    1010011101001011    1010011101001100    1010011101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42825 - 42829

  --1010011101001110    1010011101001111    1010011101010000    1010011101010001    1010011101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42830 - 42834

  --1010011101010011    1010011101010100    1010011101010101    1010011101010110    1010011101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42835 - 42839

  --1010011101011000    1010011101011001    1010011101011010    1010011101011011    1010011101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42840 - 42844

  --1010011101011101    1010011101011110    1010011101011111    1010011101100000    1010011101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42845 - 42849

  --1010011101100010    1010011101100011    1010011101100100    1010011101100101    1010011101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42850 - 42854

  --1010011101100111    1010011101101000    1010011101101001    1010011101101010    1010011101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42855 - 42859

  --1010011101101100    1010011101101101    1010011101101110    1010011101101111    1010011101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42860 - 42864

  --1010011101110001    1010011101110010    1010011101110011    1010011101110100    1010011101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42865 - 42869

  --1010011101110110    1010011101110111    1010011101111000    1010011101111001    1010011101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42870 - 42874

  --1010011101111011    1010011101111100    1010011101111101    1010011101111110    1010011101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42875 - 42879

  --1010011110000000    1010011110000001    1010011110000010    1010011110000011    1010011110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42880 - 42884

  --1010011110000101    1010011110000110    1010011110000111    1010011110001000    1010011110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42885 - 42889

  --1010011110001010    1010011110001011    1010011110001100    1010011110001101    1010011110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42890 - 42894

  --1010011110001111    1010011110010000    1010011110010001    1010011110010010    1010011110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42895 - 42899

  --1010011110010100    1010011110010101    1010011110010110    1010011110010111    1010011110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42900 - 42904

  --1010011110011001    1010011110011010    1010011110011011    1010011110011100    1010011110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42905 - 42909

  --1010011110011110    1010011110011111    1010011110100000    1010011110100001    1010011110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42910 - 42914

  --1010011110100011    1010011110100100    1010011110100101    1010011110100110    1010011110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42915 - 42919

  --1010011110101000    1010011110101001    1010011110101010    1010011110101011    1010011110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42920 - 42924

  --1010011110101101    1010011110101110    1010011110101111    1010011110110000    1010011110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42925 - 42929

  --1010011110110010    1010011110110011    1010011110110100    1010011110110101    1010011110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42930 - 42934

  --1010011110110111    1010011110111000    1010011110111001    1010011110111010    1010011110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42935 - 42939

  --1010011110111100    1010011110111101    1010011110111110    1010011110111111    1010011111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42940 - 42944

  --1010011111000001    1010011111000010    1010011111000011    1010011111000100    1010011111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42945 - 42949

  --1010011111000110    1010011111000111    1010011111001000    1010011111001001    1010011111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42950 - 42954

  --1010011111001011    1010011111001100    1010011111001101    1010011111001110    1010011111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42955 - 42959

  --1010011111010000    1010011111010001    1010011111010010    1010011111010011    1010011111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42960 - 42964

  --1010011111010101    1010011111010110    1010011111010111    1010011111011000    1010011111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42965 - 42969

  --1010011111011010    1010011111011011    1010011111011100    1010011111011101    1010011111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42970 - 42974

  --1010011111011111    1010011111100000    1010011111100001    1010011111100010    1010011111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42975 - 42979

  --1010011111100100    1010011111100101    1010011111100110    1010011111100111    1010011111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42980 - 42984

  --1010011111101001    1010011111101010    1010011111101011    1010011111101100    1010011111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42985 - 42989

  --1010011111101110    1010011111101111    1010011111110000    1010011111110001    1010011111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42990 - 42994

  --1010011111110011    1010011111110100    1010011111110101    1010011111110110    1010011111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 42995 - 42999

  --1010011111111000    1010011111111001    1010011111111010    1010011111111011    1010011111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43000 - 43004

  --1010011111111101    1010011111111110    1010011111111111    1010100000000000    1010100000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43005 - 43009

  --1010100000000010    1010100000000011    1010100000000100    1010100000000101    1010100000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43010 - 43014

  --1010100000000111    1010100000001000    1010100000001001    1010100000001010    1010100000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43015 - 43019

  --1010100000001100    1010100000001101    1010100000001110    1010100000001111    1010100000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43020 - 43024

  --1010100000010001    1010100000010010    1010100000010011    1010100000010100    1010100000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43025 - 43029

  --1010100000010110    1010100000010111    1010100000011000    1010100000011001    1010100000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43030 - 43034

  --1010100000011011    1010100000011100    1010100000011101    1010100000011110    1010100000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43035 - 43039

  --1010100000100000    1010100000100001    1010100000100010    1010100000100011    1010100000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43040 - 43044

  --1010100000100101    1010100000100110    1010100000100111    1010100000101000    1010100000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43045 - 43049

  --1010100000101010    1010100000101011    1010100000101100    1010100000101101    1010100000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43050 - 43054

  --1010100000101111    1010100000110000    1010100000110001    1010100000110010    1010100000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43055 - 43059

  --1010100000110100    1010100000110101    1010100000110110    1010100000110111    1010100000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43060 - 43064

  --1010100000111001    1010100000111010    1010100000111011    1010100000111100    1010100000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43065 - 43069

  --1010100000111110    1010100000111111    1010100001000000    1010100001000001    1010100001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43070 - 43074

  --1010100001000011    1010100001000100    1010100001000101    1010100001000110    1010100001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43075 - 43079

  --1010100001001000    1010100001001001    1010100001001010    1010100001001011    1010100001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43080 - 43084

  --1010100001001101    1010100001001110    1010100001001111    1010100001010000    1010100001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43085 - 43089

  --1010100001010010    1010100001010011    1010100001010100    1010100001010101    1010100001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43090 - 43094

  --1010100001010111    1010100001011000    1010100001011001    1010100001011010    1010100001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43095 - 43099

  --1010100001011100    1010100001011101    1010100001011110    1010100001011111    1010100001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43100 - 43104

  --1010100001100001    1010100001100010    1010100001100011    1010100001100100    1010100001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43105 - 43109

  --1010100001100110    1010100001100111    1010100001101000    1010100001101001    1010100001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43110 - 43114

  --1010100001101011    1010100001101100    1010100001101101    1010100001101110    1010100001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43115 - 43119

  --1010100001110000    1010100001110001    1010100001110010    1010100001110011    1010100001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43120 - 43124

  --1010100001110101    1010100001110110    1010100001110111    1010100001111000    1010100001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43125 - 43129

  --1010100001111010    1010100001111011    1010100001111100    1010100001111101    1010100001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43130 - 43134

  --1010100001111111    1010100010000000    1010100010000001    1010100010000010    1010100010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43135 - 43139

  --1010100010000100    1010100010000101    1010100010000110    1010100010000111    1010100010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43140 - 43144

  --1010100010001001    1010100010001010    1010100010001011    1010100010001100    1010100010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43145 - 43149

  --1010100010001110    1010100010001111    1010100010010000    1010100010010001    1010100010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43150 - 43154

  --1010100010010011    1010100010010100    1010100010010101    1010100010010110    1010100010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43155 - 43159

  --1010100010011000    1010100010011001    1010100010011010    1010100010011011    1010100010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43160 - 43164

  --1010100010011101    1010100010011110    1010100010011111    1010100010100000    1010100010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43165 - 43169

  --1010100010100010    1010100010100011    1010100010100100    1010100010100101    1010100010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43170 - 43174

  --1010100010100111    1010100010101000    1010100010101001    1010100010101010    1010100010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43175 - 43179

  --1010100010101100    1010100010101101    1010100010101110    1010100010101111    1010100010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43180 - 43184

  --1010100010110001    1010100010110010    1010100010110011    1010100010110100    1010100010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43185 - 43189

  --1010100010110110    1010100010110111    1010100010111000    1010100010111001    1010100010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43190 - 43194

  --1010100010111011    1010100010111100    1010100010111101    1010100010111110    1010100010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43195 - 43199

  --1010100011000000    1010100011000001    1010100011000010    1010100011000011    1010100011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43200 - 43204

  --1010100011000101    1010100011000110    1010100011000111    1010100011001000    1010100011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43205 - 43209

  --1010100011001010    1010100011001011    1010100011001100    1010100011001101    1010100011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43210 - 43214

  --1010100011001111    1010100011010000    1010100011010001    1010100011010010    1010100011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43215 - 43219

  --1010100011010100    1010100011010101    1010100011010110    1010100011010111    1010100011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43220 - 43224

  --1010100011011001    1010100011011010    1010100011011011    1010100011011100    1010100011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43225 - 43229

  --1010100011011110    1010100011011111    1010100011100000    1010100011100001    1010100011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43230 - 43234

  --1010100011100011    1010100011100100    1010100011100101    1010100011100110    1010100011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43235 - 43239

  --1010100011101000    1010100011101001    1010100011101010    1010100011101011    1010100011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43240 - 43244

  --1010100011101101    1010100011101110    1010100011101111    1010100011110000    1010100011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43245 - 43249

  --1010100011110010    1010100011110011    1010100011110100    1010100011110101    1010100011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43250 - 43254

  --1010100011110111    1010100011111000    1010100011111001    1010100011111010    1010100011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43255 - 43259

  --1010100011111100    1010100011111101    1010100011111110    1010100011111111    1010100100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43260 - 43264

  --1010100100000001    1010100100000010    1010100100000011    1010100100000100    1010100100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43265 - 43269

  --1010100100000110    1010100100000111    1010100100001000    1010100100001001    1010100100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43270 - 43274

  --1010100100001011    1010100100001100    1010100100001101    1010100100001110    1010100100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43275 - 43279

  --1010100100010000    1010100100010001    1010100100010010    1010100100010011    1010100100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43280 - 43284

  --1010100100010101    1010100100010110    1010100100010111    1010100100011000    1010100100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43285 - 43289

  --1010100100011010    1010100100011011    1010100100011100    1010100100011101    1010100100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43290 - 43294

  --1010100100011111    1010100100100000    1010100100100001    1010100100100010    1010100100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43295 - 43299

  --1010100100100100    1010100100100101    1010100100100110    1010100100100111    1010100100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43300 - 43304

  --1010100100101001    1010100100101010    1010100100101011    1010100100101100    1010100100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43305 - 43309

  --1010100100101110    1010100100101111    1010100100110000    1010100100110001    1010100100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43310 - 43314

  --1010100100110011    1010100100110100    1010100100110101    1010100100110110    1010100100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43315 - 43319

  --1010100100111000    1010100100111001    1010100100111010    1010100100111011    1010100100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43320 - 43324

  --1010100100111101    1010100100111110    1010100100111111    1010100101000000    1010100101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43325 - 43329

  --1010100101000010    1010100101000011    1010100101000100    1010100101000101    1010100101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43330 - 43334

  --1010100101000111    1010100101001000    1010100101001001    1010100101001010    1010100101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43335 - 43339

  --1010100101001100    1010100101001101    1010100101001110    1010100101001111    1010100101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43340 - 43344

  --1010100101010001    1010100101010010    1010100101010011    1010100101010100    1010100101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43345 - 43349

  --1010100101010110    1010100101010111    1010100101011000    1010100101011001    1010100101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43350 - 43354

  --1010100101011011    1010100101011100    1010100101011101    1010100101011110    1010100101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43355 - 43359

  --1010100101100000    1010100101100001    1010100101100010    1010100101100011    1010100101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43360 - 43364

  --1010100101100101    1010100101100110    1010100101100111    1010100101101000    1010100101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43365 - 43369

  --1010100101101010    1010100101101011    1010100101101100    1010100101101101    1010100101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43370 - 43374

  --1010100101101111    1010100101110000    1010100101110001    1010100101110010    1010100101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43375 - 43379

  --1010100101110100    1010100101110101    1010100101110110    1010100101110111    1010100101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43380 - 43384

  --1010100101111001    1010100101111010    1010100101111011    1010100101111100    1010100101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43385 - 43389

  --1010100101111110    1010100101111111    1010100110000000    1010100110000001    1010100110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43390 - 43394

  --1010100110000011    1010100110000100    1010100110000101    1010100110000110    1010100110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43395 - 43399

  --1010100110001000    1010100110001001    1010100110001010    1010100110001011    1010100110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43400 - 43404

  --1010100110001101    1010100110001110    1010100110001111    1010100110010000    1010100110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43405 - 43409

  --1010100110010010    1010100110010011    1010100110010100    1010100110010101    1010100110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43410 - 43414

  --1010100110010111    1010100110011000    1010100110011001    1010100110011010    1010100110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43415 - 43419

  --1010100110011100    1010100110011101    1010100110011110    1010100110011111    1010100110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43420 - 43424

  --1010100110100001    1010100110100010    1010100110100011    1010100110100100    1010100110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43425 - 43429

  --1010100110100110    1010100110100111    1010100110101000    1010100110101001    1010100110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43430 - 43434

  --1010100110101011    1010100110101100    1010100110101101    1010100110101110    1010100110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43435 - 43439

  --1010100110110000    1010100110110001    1010100110110010    1010100110110011    1010100110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43440 - 43444

  --1010100110110101    1010100110110110    1010100110110111    1010100110111000    1010100110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43445 - 43449

  --1010100110111010    1010100110111011    1010100110111100    1010100110111101    1010100110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43450 - 43454

  --1010100110111111    1010100111000000    1010100111000001    1010100111000010    1010100111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43455 - 43459

  --1010100111000100    1010100111000101    1010100111000110    1010100111000111    1010100111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43460 - 43464

  --1010100111001001    1010100111001010    1010100111001011    1010100111001100    1010100111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43465 - 43469

  --1010100111001110    1010100111001111    1010100111010000    1010100111010001    1010100111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43470 - 43474

  --1010100111010011    1010100111010100    1010100111010101    1010100111010110    1010100111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43475 - 43479

  --1010100111011000    1010100111011001    1010100111011010    1010100111011011    1010100111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43480 - 43484

  --1010100111011101    1010100111011110    1010100111011111    1010100111100000    1010100111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43485 - 43489

  --1010100111100010    1010100111100011    1010100111100100    1010100111100101    1010100111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43490 - 43494

  --1010100111100111    1010100111101000    1010100111101001    1010100111101010    1010100111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43495 - 43499

  --1010100111101100    1010100111101101    1010100111101110    1010100111101111    1010100111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43500 - 43504

  --1010100111110001    1010100111110010    1010100111110011    1010100111110100    1010100111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43505 - 43509

  --1010100111110110    1010100111110111    1010100111111000    1010100111111001    1010100111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43510 - 43514

  --1010100111111011    1010100111111100    1010100111111101    1010100111111110    1010100111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43515 - 43519

  --1010101000000000    1010101000000001    1010101000000010    1010101000000011    1010101000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43520 - 43524

  --1010101000000101    1010101000000110    1010101000000111    1010101000001000    1010101000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43525 - 43529

  --1010101000001010    1010101000001011    1010101000001100    1010101000001101    1010101000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43530 - 43534

  --1010101000001111    1010101000010000    1010101000010001    1010101000010010    1010101000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43535 - 43539

  --1010101000010100    1010101000010101    1010101000010110    1010101000010111    1010101000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43540 - 43544

  --1010101000011001    1010101000011010    1010101000011011    1010101000011100    1010101000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43545 - 43549

  --1010101000011110    1010101000011111    1010101000100000    1010101000100001    1010101000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43550 - 43554

  --1010101000100011    1010101000100100    1010101000100101    1010101000100110    1010101000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43555 - 43559

  --1010101000101000    1010101000101001    1010101000101010    1010101000101011    1010101000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43560 - 43564

  --1010101000101101    1010101000101110    1010101000101111    1010101000110000    1010101000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43565 - 43569

  --1010101000110010    1010101000110011    1010101000110100    1010101000110101    1010101000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43570 - 43574

  --1010101000110111    1010101000111000    1010101000111001    1010101000111010    1010101000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43575 - 43579

  --1010101000111100    1010101000111101    1010101000111110    1010101000111111    1010101001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43580 - 43584

  --1010101001000001    1010101001000010    1010101001000011    1010101001000100    1010101001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43585 - 43589

  --1010101001000110    1010101001000111    1010101001001000    1010101001001001    1010101001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43590 - 43594

  --1010101001001011    1010101001001100    1010101001001101    1010101001001110    1010101001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43595 - 43599

  --1010101001010000    1010101001010001    1010101001010010    1010101001010011    1010101001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43600 - 43604

  --1010101001010101    1010101001010110    1010101001010111    1010101001011000    1010101001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43605 - 43609

  --1010101001011010    1010101001011011    1010101001011100    1010101001011101    1010101001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43610 - 43614

  --1010101001011111    1010101001100000    1010101001100001    1010101001100010    1010101001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43615 - 43619

  --1010101001100100    1010101001100101    1010101001100110    1010101001100111    1010101001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43620 - 43624

  --1010101001101001    1010101001101010    1010101001101011    1010101001101100    1010101001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43625 - 43629

  --1010101001101110    1010101001101111    1010101001110000    1010101001110001    1010101001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43630 - 43634

  --1010101001110011    1010101001110100    1010101001110101    1010101001110110    1010101001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43635 - 43639

  --1010101001111000    1010101001111001    1010101001111010    1010101001111011    1010101001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43640 - 43644

  --1010101001111101    1010101001111110    1010101001111111    1010101010000000    1010101010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43645 - 43649

  --1010101010000010    1010101010000011    1010101010000100    1010101010000101    1010101010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43650 - 43654

  --1010101010000111    1010101010001000    1010101010001001    1010101010001010    1010101010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43655 - 43659

  --1010101010001100    1010101010001101    1010101010001110    1010101010001111    1010101010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43660 - 43664

  --1010101010010001    1010101010010010    1010101010010011    1010101010010100    1010101010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43665 - 43669

  --1010101010010110    1010101010010111    1010101010011000    1010101010011001    1010101010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43670 - 43674

  --1010101010011011    1010101010011100    1010101010011101    1010101010011110    1010101010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43675 - 43679

  --1010101010100000    1010101010100001    1010101010100010    1010101010100011    1010101010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43680 - 43684

  --1010101010100101    1010101010100110    1010101010100111    1010101010101000    1010101010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43685 - 43689

  --1010101010101010    1010101010101011    1010101010101100    1010101010101101    1010101010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43690 - 43694

  --1010101010101111    1010101010110000    1010101010110001    1010101010110010    1010101010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43695 - 43699

  --1010101010110100    1010101010110101    1010101010110110    1010101010110111    1010101010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43700 - 43704

  --1010101010111001    1010101010111010    1010101010111011    1010101010111100    1010101010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43705 - 43709

  --1010101010111110    1010101010111111    1010101011000000    1010101011000001    1010101011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43710 - 43714

  --1010101011000011    1010101011000100    1010101011000101    1010101011000110    1010101011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43715 - 43719

  --1010101011001000    1010101011001001    1010101011001010    1010101011001011    1010101011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43720 - 43724

  --1010101011001101    1010101011001110    1010101011001111    1010101011010000    1010101011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43725 - 43729

  --1010101011010010    1010101011010011    1010101011010100    1010101011010101    1010101011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43730 - 43734

  --1010101011010111    1010101011011000    1010101011011001    1010101011011010    1010101011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43735 - 43739

  --1010101011011100    1010101011011101    1010101011011110    1010101011011111    1010101011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43740 - 43744

  --1010101011100001    1010101011100010    1010101011100011    1010101011100100    1010101011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43745 - 43749

  --1010101011100110    1010101011100111    1010101011101000    1010101011101001    1010101011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43750 - 43754

  --1010101011101011    1010101011101100    1010101011101101    1010101011101110    1010101011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43755 - 43759

  --1010101011110000    1010101011110001    1010101011110010    1010101011110011    1010101011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43760 - 43764

  --1010101011110101    1010101011110110    1010101011110111    1010101011111000    1010101011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43765 - 43769

  --1010101011111010    1010101011111011    1010101011111100    1010101011111101    1010101011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43770 - 43774

  --1010101011111111    1010101100000000    1010101100000001    1010101100000010    1010101100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43775 - 43779

  --1010101100000100    1010101100000101    1010101100000110    1010101100000111    1010101100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43780 - 43784

  --1010101100001001    1010101100001010    1010101100001011    1010101100001100    1010101100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43785 - 43789

  --1010101100001110    1010101100001111    1010101100010000    1010101100010001    1010101100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43790 - 43794

  --1010101100010011    1010101100010100    1010101100010101    1010101100010110    1010101100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43795 - 43799

  --1010101100011000    1010101100011001    1010101100011010    1010101100011011    1010101100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43800 - 43804

  --1010101100011101    1010101100011110    1010101100011111    1010101100100000    1010101100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43805 - 43809

  --1010101100100010    1010101100100011    1010101100100100    1010101100100101    1010101100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43810 - 43814

  --1010101100100111    1010101100101000    1010101100101001    1010101100101010    1010101100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43815 - 43819

  --1010101100101100    1010101100101101    1010101100101110    1010101100101111    1010101100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43820 - 43824

  --1010101100110001    1010101100110010    1010101100110011    1010101100110100    1010101100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43825 - 43829

  --1010101100110110    1010101100110111    1010101100111000    1010101100111001    1010101100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43830 - 43834

  --1010101100111011    1010101100111100    1010101100111101    1010101100111110    1010101100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43835 - 43839

  --1010101101000000    1010101101000001    1010101101000010    1010101101000011    1010101101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43840 - 43844

  --1010101101000101    1010101101000110    1010101101000111    1010101101001000    1010101101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43845 - 43849

  --1010101101001010    1010101101001011    1010101101001100    1010101101001101    1010101101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43850 - 43854

  --1010101101001111    1010101101010000    1010101101010001    1010101101010010    1010101101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43855 - 43859

  --1010101101010100    1010101101010101    1010101101010110    1010101101010111    1010101101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43860 - 43864

  --1010101101011001    1010101101011010    1010101101011011    1010101101011100    1010101101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43865 - 43869

  --1010101101011110    1010101101011111    1010101101100000    1010101101100001    1010101101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43870 - 43874

  --1010101101100011    1010101101100100    1010101101100101    1010101101100110    1010101101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43875 - 43879

  --1010101101101000    1010101101101001    1010101101101010    1010101101101011    1010101101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43880 - 43884

  --1010101101101101    1010101101101110    1010101101101111    1010101101110000    1010101101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43885 - 43889

  --1010101101110010    1010101101110011    1010101101110100    1010101101110101    1010101101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43890 - 43894

  --1010101101110111    1010101101111000    1010101101111001    1010101101111010    1010101101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43895 - 43899

  --1010101101111100    1010101101111101    1010101101111110    1010101101111111    1010101110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43900 - 43904

  --1010101110000001    1010101110000010    1010101110000011    1010101110000100    1010101110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43905 - 43909

  --1010101110000110    1010101110000111    1010101110001000    1010101110001001    1010101110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43910 - 43914

  --1010101110001011    1010101110001100    1010101110001101    1010101110001110    1010101110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43915 - 43919

  --1010101110010000    1010101110010001    1010101110010010    1010101110010011    1010101110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43920 - 43924

  --1010101110010101    1010101110010110    1010101110010111    1010101110011000    1010101110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43925 - 43929

  --1010101110011010    1010101110011011    1010101110011100    1010101110011101    1010101110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43930 - 43934

  --1010101110011111    1010101110100000    1010101110100001    1010101110100010    1010101110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43935 - 43939

  --1010101110100100    1010101110100101    1010101110100110    1010101110100111    1010101110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43940 - 43944

  --1010101110101001    1010101110101010    1010101110101011    1010101110101100    1010101110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43945 - 43949

  --1010101110101110    1010101110101111    1010101110110000    1010101110110001    1010101110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43950 - 43954

  --1010101110110011    1010101110110100    1010101110110101    1010101110110110    1010101110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43955 - 43959

  --1010101110111000    1010101110111001    1010101110111010    1010101110111011    1010101110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43960 - 43964

  --1010101110111101    1010101110111110    1010101110111111    1010101111000000    1010101111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43965 - 43969

  --1010101111000010    1010101111000011    1010101111000100    1010101111000101    1010101111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43970 - 43974

  --1010101111000111    1010101111001000    1010101111001001    1010101111001010    1010101111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43975 - 43979

  --1010101111001100    1010101111001101    1010101111001110    1010101111001111    1010101111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43980 - 43984

  --1010101111010001    1010101111010010    1010101111010011    1010101111010100    1010101111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43985 - 43989

  --1010101111010110    1010101111010111    1010101111011000    1010101111011001    1010101111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43990 - 43994

  --1010101111011011    1010101111011100    1010101111011101    1010101111011110    1010101111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 43995 - 43999

  --1010101111100000    1010101111100001    1010101111100010    1010101111100011    1010101111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44000 - 44004

  --1010101111100101    1010101111100110    1010101111100111    1010101111101000    1010101111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44005 - 44009

  --1010101111101010    1010101111101011    1010101111101100    1010101111101101    1010101111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44010 - 44014

  --1010101111101111    1010101111110000    1010101111110001    1010101111110010    1010101111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44015 - 44019

  --1010101111110100    1010101111110101    1010101111110110    1010101111110111    1010101111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44020 - 44024

  --1010101111111001    1010101111111010    1010101111111011    1010101111111100    1010101111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44025 - 44029

  --1010101111111110    1010101111111111    1010110000000000    1010110000000001    1010110000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44030 - 44034

  --1010110000000011    1010110000000100    1010110000000101    1010110000000110    1010110000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44035 - 44039

  --1010110000001000    1010110000001001    1010110000001010    1010110000001011    1010110000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44040 - 44044

  --1010110000001101    1010110000001110    1010110000001111    1010110000010000    1010110000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44045 - 44049

  --1010110000010010    1010110000010011    1010110000010100    1010110000010101    1010110000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44050 - 44054

  --1010110000010111    1010110000011000    1010110000011001    1010110000011010    1010110000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44055 - 44059

  --1010110000011100    1010110000011101    1010110000011110    1010110000011111    1010110000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44060 - 44064

  --1010110000100001    1010110000100010    1010110000100011    1010110000100100    1010110000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44065 - 44069

  --1010110000100110    1010110000100111    1010110000101000    1010110000101001    1010110000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44070 - 44074

  --1010110000101011    1010110000101100    1010110000101101    1010110000101110    1010110000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44075 - 44079

  --1010110000110000    1010110000110001    1010110000110010    1010110000110011    1010110000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44080 - 44084

  --1010110000110101    1010110000110110    1010110000110111    1010110000111000    1010110000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44085 - 44089

  --1010110000111010    1010110000111011    1010110000111100    1010110000111101    1010110000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44090 - 44094

  --1010110000111111    1010110001000000    1010110001000001    1010110001000010    1010110001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44095 - 44099

  --1010110001000100    1010110001000101    1010110001000110    1010110001000111    1010110001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44100 - 44104

  --1010110001001001    1010110001001010    1010110001001011    1010110001001100    1010110001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44105 - 44109

  --1010110001001110    1010110001001111    1010110001010000    1010110001010001    1010110001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44110 - 44114

  --1010110001010011    1010110001010100    1010110001010101    1010110001010110    1010110001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44115 - 44119

  --1010110001011000    1010110001011001    1010110001011010    1010110001011011    1010110001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44120 - 44124

  --1010110001011101    1010110001011110    1010110001011111    1010110001100000    1010110001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44125 - 44129

  --1010110001100010    1010110001100011    1010110001100100    1010110001100101    1010110001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44130 - 44134

  --1010110001100111    1010110001101000    1010110001101001    1010110001101010    1010110001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44135 - 44139

  --1010110001101100    1010110001101101    1010110001101110    1010110001101111    1010110001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44140 - 44144

  --1010110001110001    1010110001110010    1010110001110011    1010110001110100    1010110001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44145 - 44149

  --1010110001110110    1010110001110111    1010110001111000    1010110001111001    1010110001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44150 - 44154

  --1010110001111011    1010110001111100    1010110001111101    1010110001111110    1010110001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44155 - 44159

  --1010110010000000    1010110010000001    1010110010000010    1010110010000011    1010110010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44160 - 44164

  --1010110010000101    1010110010000110    1010110010000111    1010110010001000    1010110010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44165 - 44169

  --1010110010001010    1010110010001011    1010110010001100    1010110010001101    1010110010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44170 - 44174

  --1010110010001111    1010110010010000    1010110010010001    1010110010010010    1010110010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44175 - 44179

  --1010110010010100    1010110010010101    1010110010010110    1010110010010111    1010110010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44180 - 44184

  --1010110010011001    1010110010011010    1010110010011011    1010110010011100    1010110010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44185 - 44189

  --1010110010011110    1010110010011111    1010110010100000    1010110010100001    1010110010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44190 - 44194

  --1010110010100011    1010110010100100    1010110010100101    1010110010100110    1010110010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44195 - 44199

  --1010110010101000    1010110010101001    1010110010101010    1010110010101011    1010110010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44200 - 44204

  --1010110010101101    1010110010101110    1010110010101111    1010110010110000    1010110010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44205 - 44209

  --1010110010110010    1010110010110011    1010110010110100    1010110010110101    1010110010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44210 - 44214

  --1010110010110111    1010110010111000    1010110010111001    1010110010111010    1010110010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44215 - 44219

  --1010110010111100    1010110010111101    1010110010111110    1010110010111111    1010110011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44220 - 44224

  --1010110011000001    1010110011000010    1010110011000011    1010110011000100    1010110011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44225 - 44229

  --1010110011000110    1010110011000111    1010110011001000    1010110011001001    1010110011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44230 - 44234

  --1010110011001011    1010110011001100    1010110011001101    1010110011001110    1010110011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44235 - 44239

  --1010110011010000    1010110011010001    1010110011010010    1010110011010011    1010110011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44240 - 44244

  --1010110011010101    1010110011010110    1010110011010111    1010110011011000    1010110011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44245 - 44249

  --1010110011011010    1010110011011011    1010110011011100    1010110011011101    1010110011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44250 - 44254

  --1010110011011111    1010110011100000    1010110011100001    1010110011100010    1010110011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44255 - 44259

  --1010110011100100    1010110011100101    1010110011100110    1010110011100111    1010110011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44260 - 44264

  --1010110011101001    1010110011101010    1010110011101011    1010110011101100    1010110011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44265 - 44269

  --1010110011101110    1010110011101111    1010110011110000    1010110011110001    1010110011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44270 - 44274

  --1010110011110011    1010110011110100    1010110011110101    1010110011110110    1010110011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44275 - 44279

  --1010110011111000    1010110011111001    1010110011111010    1010110011111011    1010110011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44280 - 44284

  --1010110011111101    1010110011111110    1010110011111111    1010110100000000    1010110100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44285 - 44289

  --1010110100000010    1010110100000011    1010110100000100    1010110100000101    1010110100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44290 - 44294

  --1010110100000111    1010110100001000    1010110100001001    1010110100001010    1010110100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44295 - 44299

  --1010110100001100    1010110100001101    1010110100001110    1010110100001111    1010110100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44300 - 44304

  --1010110100010001    1010110100010010    1010110100010011    1010110100010100    1010110100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44305 - 44309

  --1010110100010110    1010110100010111    1010110100011000    1010110100011001    1010110100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44310 - 44314

  --1010110100011011    1010110100011100    1010110100011101    1010110100011110    1010110100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44315 - 44319

  --1010110100100000    1010110100100001    1010110100100010    1010110100100011    1010110100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44320 - 44324

  --1010110100100101    1010110100100110    1010110100100111    1010110100101000    1010110100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44325 - 44329

  --1010110100101010    1010110100101011    1010110100101100    1010110100101101    1010110100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44330 - 44334

  --1010110100101111    1010110100110000    1010110100110001    1010110100110010    1010110100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44335 - 44339

  --1010110100110100    1010110100110101    1010110100110110    1010110100110111    1010110100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44340 - 44344

  --1010110100111001    1010110100111010    1010110100111011    1010110100111100    1010110100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44345 - 44349

  --1010110100111110    1010110100111111    1010110101000000    1010110101000001    1010110101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44350 - 44354

  --1010110101000011    1010110101000100    1010110101000101    1010110101000110    1010110101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44355 - 44359

  --1010110101001000    1010110101001001    1010110101001010    1010110101001011    1010110101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44360 - 44364

  --1010110101001101    1010110101001110    1010110101001111    1010110101010000    1010110101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44365 - 44369

  --1010110101010010    1010110101010011    1010110101010100    1010110101010101    1010110101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44370 - 44374

  --1010110101010111    1010110101011000    1010110101011001    1010110101011010    1010110101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44375 - 44379

  --1010110101011100    1010110101011101    1010110101011110    1010110101011111    1010110101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44380 - 44384

  --1010110101100001    1010110101100010    1010110101100011    1010110101100100    1010110101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44385 - 44389

  --1010110101100110    1010110101100111    1010110101101000    1010110101101001    1010110101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44390 - 44394

  --1010110101101011    1010110101101100    1010110101101101    1010110101101110    1010110101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44395 - 44399

  --1010110101110000    1010110101110001    1010110101110010    1010110101110011    1010110101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44400 - 44404

  --1010110101110101    1010110101110110    1010110101110111    1010110101111000    1010110101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44405 - 44409

  --1010110101111010    1010110101111011    1010110101111100    1010110101111101    1010110101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44410 - 44414

  --1010110101111111    1010110110000000    1010110110000001    1010110110000010    1010110110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44415 - 44419

  --1010110110000100    1010110110000101    1010110110000110    1010110110000111    1010110110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44420 - 44424

  --1010110110001001    1010110110001010    1010110110001011    1010110110001100    1010110110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44425 - 44429

  --1010110110001110    1010110110001111    1010110110010000    1010110110010001    1010110110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44430 - 44434

  --1010110110010011    1010110110010100    1010110110010101    1010110110010110    1010110110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44435 - 44439

  --1010110110011000    1010110110011001    1010110110011010    1010110110011011    1010110110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44440 - 44444

  --1010110110011101    1010110110011110    1010110110011111    1010110110100000    1010110110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44445 - 44449

  --1010110110100010    1010110110100011    1010110110100100    1010110110100101    1010110110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44450 - 44454

  --1010110110100111    1010110110101000    1010110110101001    1010110110101010    1010110110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44455 - 44459

  --1010110110101100    1010110110101101    1010110110101110    1010110110101111    1010110110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44460 - 44464

  --1010110110110001    1010110110110010    1010110110110011    1010110110110100    1010110110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44465 - 44469

  --1010110110110110    1010110110110111    1010110110111000    1010110110111001    1010110110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44470 - 44474

  --1010110110111011    1010110110111100    1010110110111101    1010110110111110    1010110110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44475 - 44479

  --1010110111000000    1010110111000001    1010110111000010    1010110111000011    1010110111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44480 - 44484

  --1010110111000101    1010110111000110    1010110111000111    1010110111001000    1010110111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44485 - 44489

  --1010110111001010    1010110111001011    1010110111001100    1010110111001101    1010110111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44490 - 44494

  --1010110111001111    1010110111010000    1010110111010001    1010110111010010    1010110111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44495 - 44499

  --1010110111010100    1010110111010101    1010110111010110    1010110111010111    1010110111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44500 - 44504

  --1010110111011001    1010110111011010    1010110111011011    1010110111011100    1010110111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44505 - 44509

  --1010110111011110    1010110111011111    1010110111100000    1010110111100001    1010110111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44510 - 44514

  --1010110111100011    1010110111100100    1010110111100101    1010110111100110    1010110111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44515 - 44519

  --1010110111101000    1010110111101001    1010110111101010    1010110111101011    1010110111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44520 - 44524

  --1010110111101101    1010110111101110    1010110111101111    1010110111110000    1010110111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44525 - 44529

  --1010110111110010    1010110111110011    1010110111110100    1010110111110101    1010110111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44530 - 44534

  --1010110111110111    1010110111111000    1010110111111001    1010110111111010    1010110111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44535 - 44539

  --1010110111111100    1010110111111101    1010110111111110    1010110111111111    1010111000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44540 - 44544

  --1010111000000001    1010111000000010    1010111000000011    1010111000000100    1010111000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44545 - 44549

  --1010111000000110    1010111000000111    1010111000001000    1010111000001001    1010111000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44550 - 44554

  --1010111000001011    1010111000001100    1010111000001101    1010111000001110    1010111000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44555 - 44559

  --1010111000010000    1010111000010001    1010111000010010    1010111000010011    1010111000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44560 - 44564

  --1010111000010101    1010111000010110    1010111000010111    1010111000011000    1010111000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44565 - 44569

  --1010111000011010    1010111000011011    1010111000011100    1010111000011101    1010111000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44570 - 44574

  --1010111000011111    1010111000100000    1010111000100001    1010111000100010    1010111000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44575 - 44579

  --1010111000100100    1010111000100101    1010111000100110    1010111000100111    1010111000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44580 - 44584

  --1010111000101001    1010111000101010    1010111000101011    1010111000101100    1010111000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44585 - 44589

  --1010111000101110    1010111000101111    1010111000110000    1010111000110001    1010111000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44590 - 44594

  --1010111000110011    1010111000110100    1010111000110101    1010111000110110    1010111000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44595 - 44599

  --1010111000111000    1010111000111001    1010111000111010    1010111000111011    1010111000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44600 - 44604

  --1010111000111101    1010111000111110    1010111000111111    1010111001000000    1010111001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44605 - 44609

  --1010111001000010    1010111001000011    1010111001000100    1010111001000101    1010111001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44610 - 44614

  --1010111001000111    1010111001001000    1010111001001001    1010111001001010    1010111001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44615 - 44619

  --1010111001001100    1010111001001101    1010111001001110    1010111001001111    1010111001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44620 - 44624

  --1010111001010001    1010111001010010    1010111001010011    1010111001010100    1010111001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44625 - 44629

  --1010111001010110    1010111001010111    1010111001011000    1010111001011001    1010111001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44630 - 44634

  --1010111001011011    1010111001011100    1010111001011101    1010111001011110    1010111001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44635 - 44639

  --1010111001100000    1010111001100001    1010111001100010    1010111001100011    1010111001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44640 - 44644

  --1010111001100101    1010111001100110    1010111001100111    1010111001101000    1010111001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44645 - 44649

  --1010111001101010    1010111001101011    1010111001101100    1010111001101101    1010111001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44650 - 44654

  --1010111001101111    1010111001110000    1010111001110001    1010111001110010    1010111001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44655 - 44659

  --1010111001110100    1010111001110101    1010111001110110    1010111001110111    1010111001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44660 - 44664

  --1010111001111001    1010111001111010    1010111001111011    1010111001111100    1010111001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44665 - 44669

  --1010111001111110    1010111001111111    1010111010000000    1010111010000001    1010111010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44670 - 44674

  --1010111010000011    1010111010000100    1010111010000101    1010111010000110    1010111010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44675 - 44679

  --1010111010001000    1010111010001001    1010111010001010    1010111010001011    1010111010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44680 - 44684

  --1010111010001101    1010111010001110    1010111010001111    1010111010010000    1010111010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44685 - 44689

  --1010111010010010    1010111010010011    1010111010010100    1010111010010101    1010111010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44690 - 44694

  --1010111010010111    1010111010011000    1010111010011001    1010111010011010    1010111010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44695 - 44699

  --1010111010011100    1010111010011101    1010111010011110    1010111010011111    1010111010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44700 - 44704

  --1010111010100001    1010111010100010    1010111010100011    1010111010100100    1010111010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44705 - 44709

  --1010111010100110    1010111010100111    1010111010101000    1010111010101001    1010111010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44710 - 44714

  --1010111010101011    1010111010101100    1010111010101101    1010111010101110    1010111010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44715 - 44719

  --1010111010110000    1010111010110001    1010111010110010    1010111010110011    1010111010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44720 - 44724

  --1010111010110101    1010111010110110    1010111010110111    1010111010111000    1010111010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44725 - 44729

  --1010111010111010    1010111010111011    1010111010111100    1010111010111101    1010111010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44730 - 44734

  --1010111010111111    1010111011000000    1010111011000001    1010111011000010    1010111011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44735 - 44739

  --1010111011000100    1010111011000101    1010111011000110    1010111011000111    1010111011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44740 - 44744

  --1010111011001001    1010111011001010    1010111011001011    1010111011001100    1010111011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44745 - 44749

  --1010111011001110    1010111011001111    1010111011010000    1010111011010001    1010111011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44750 - 44754

  --1010111011010011    1010111011010100    1010111011010101    1010111011010110    1010111011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44755 - 44759

  --1010111011011000    1010111011011001    1010111011011010    1010111011011011    1010111011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44760 - 44764

  --1010111011011101    1010111011011110    1010111011011111    1010111011100000    1010111011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44765 - 44769

  --1010111011100010    1010111011100011    1010111011100100    1010111011100101    1010111011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44770 - 44774

  --1010111011100111    1010111011101000    1010111011101001    1010111011101010    1010111011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44775 - 44779

  --1010111011101100    1010111011101101    1010111011101110    1010111011101111    1010111011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44780 - 44784

  --1010111011110001    1010111011110010    1010111011110011    1010111011110100    1010111011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44785 - 44789

  --1010111011110110    1010111011110111    1010111011111000    1010111011111001    1010111011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44790 - 44794

  --1010111011111011    1010111011111100    1010111011111101    1010111011111110    1010111011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44795 - 44799

  --1010111100000000    1010111100000001    1010111100000010    1010111100000011    1010111100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44800 - 44804

  --1010111100000101    1010111100000110    1010111100000111    1010111100001000    1010111100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44805 - 44809

  --1010111100001010    1010111100001011    1010111100001100    1010111100001101    1010111100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44810 - 44814

  --1010111100001111    1010111100010000    1010111100010001    1010111100010010    1010111100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44815 - 44819

  --1010111100010100    1010111100010101    1010111100010110    1010111100010111    1010111100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44820 - 44824

  --1010111100011001    1010111100011010    1010111100011011    1010111100011100    1010111100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44825 - 44829

  --1010111100011110    1010111100011111    1010111100100000    1010111100100001    1010111100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44830 - 44834

  --1010111100100011    1010111100100100    1010111100100101    1010111100100110    1010111100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44835 - 44839

  --1010111100101000    1010111100101001    1010111100101010    1010111100101011    1010111100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44840 - 44844

  --1010111100101101    1010111100101110    1010111100101111    1010111100110000    1010111100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44845 - 44849

  --1010111100110010    1010111100110011    1010111100110100    1010111100110101    1010111100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44850 - 44854

  --1010111100110111    1010111100111000    1010111100111001    1010111100111010    1010111100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44855 - 44859

  --1010111100111100    1010111100111101    1010111100111110    1010111100111111    1010111101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44860 - 44864

  --1010111101000001    1010111101000010    1010111101000011    1010111101000100    1010111101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44865 - 44869

  --1010111101000110    1010111101000111    1010111101001000    1010111101001001    1010111101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44870 - 44874

  --1010111101001011    1010111101001100    1010111101001101    1010111101001110    1010111101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44875 - 44879

  --1010111101010000    1010111101010001    1010111101010010    1010111101010011    1010111101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44880 - 44884

  --1010111101010101    1010111101010110    1010111101010111    1010111101011000    1010111101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44885 - 44889

  --1010111101011010    1010111101011011    1010111101011100    1010111101011101    1010111101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44890 - 44894

  --1010111101011111    1010111101100000    1010111101100001    1010111101100010    1010111101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44895 - 44899

  --1010111101100100    1010111101100101    1010111101100110    1010111101100111    1010111101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44900 - 44904

  --1010111101101001    1010111101101010    1010111101101011    1010111101101100    1010111101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44905 - 44909

  --1010111101101110    1010111101101111    1010111101110000    1010111101110001    1010111101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44910 - 44914

  --1010111101110011    1010111101110100    1010111101110101    1010111101110110    1010111101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44915 - 44919

  --1010111101111000    1010111101111001    1010111101111010    1010111101111011    1010111101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44920 - 44924

  --1010111101111101    1010111101111110    1010111101111111    1010111110000000    1010111110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44925 - 44929

  --1010111110000010    1010111110000011    1010111110000100    1010111110000101    1010111110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44930 - 44934

  --1010111110000111    1010111110001000    1010111110001001    1010111110001010    1010111110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44935 - 44939

  --1010111110001100    1010111110001101    1010111110001110    1010111110001111    1010111110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44940 - 44944

  --1010111110010001    1010111110010010    1010111110010011    1010111110010100    1010111110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44945 - 44949

  --1010111110010110    1010111110010111    1010111110011000    1010111110011001    1010111110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44950 - 44954

  --1010111110011011    1010111110011100    1010111110011101    1010111110011110    1010111110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44955 - 44959

  --1010111110100000    1010111110100001    1010111110100010    1010111110100011    1010111110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44960 - 44964

  --1010111110100101    1010111110100110    1010111110100111    1010111110101000    1010111110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44965 - 44969

  --1010111110101010    1010111110101011    1010111110101100    1010111110101101    1010111110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44970 - 44974

  --1010111110101111    1010111110110000    1010111110110001    1010111110110010    1010111110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44975 - 44979

  --1010111110110100    1010111110110101    1010111110110110    1010111110110111    1010111110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44980 - 44984

  --1010111110111001    1010111110111010    1010111110111011    1010111110111100    1010111110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44985 - 44989

  --1010111110111110    1010111110111111    1010111111000000    1010111111000001    1010111111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44990 - 44994

  --1010111111000011    1010111111000100    1010111111000101    1010111111000110    1010111111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 44995 - 44999

  --1010111111001000    1010111111001001    1010111111001010    1010111111001011    1010111111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45000 - 45004

  --1010111111001101    1010111111001110    1010111111001111    1010111111010000    1010111111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45005 - 45009

  --1010111111010010    1010111111010011    1010111111010100    1010111111010101    1010111111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45010 - 45014

  --1010111111010111    1010111111011000    1010111111011001    1010111111011010    1010111111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45015 - 45019

  --1010111111011100    1010111111011101    1010111111011110    1010111111011111    1010111111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45020 - 45024

  --1010111111100001    1010111111100010    1010111111100011    1010111111100100    1010111111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45025 - 45029

  --1010111111100110    1010111111100111    1010111111101000    1010111111101001    1010111111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45030 - 45034

  --1010111111101011    1010111111101100    1010111111101101    1010111111101110    1010111111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45035 - 45039

  --1010111111110000    1010111111110001    1010111111110010    1010111111110011    1010111111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45040 - 45044

  --1010111111110101    1010111111110110    1010111111110111    1010111111111000    1010111111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45045 - 45049

  --1010111111111010    1010111111111011    1010111111111100    1010111111111101    1010111111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45050 - 45054

  --1010111111111111    1011000000000000    1011000000000001    1011000000000010    1011000000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45055 - 45059

  --1011000000000100    1011000000000101    1011000000000110    1011000000000111    1011000000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45060 - 45064

  --1011000000001001    1011000000001010    1011000000001011    1011000000001100    1011000000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45065 - 45069

  --1011000000001110    1011000000001111    1011000000010000    1011000000010001    1011000000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45070 - 45074

  --1011000000010011    1011000000010100    1011000000010101    1011000000010110    1011000000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45075 - 45079

  --1011000000011000    1011000000011001    1011000000011010    1011000000011011    1011000000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45080 - 45084

  --1011000000011101    1011000000011110    1011000000011111    1011000000100000    1011000000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45085 - 45089

  --1011000000100010    1011000000100011    1011000000100100    1011000000100101    1011000000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45090 - 45094

  --1011000000100111    1011000000101000    1011000000101001    1011000000101010    1011000000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45095 - 45099

  --1011000000101100    1011000000101101    1011000000101110    1011000000101111    1011000000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45100 - 45104

  --1011000000110001    1011000000110010    1011000000110011    1011000000110100    1011000000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45105 - 45109

  --1011000000110110    1011000000110111    1011000000111000    1011000000111001    1011000000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45110 - 45114

  --1011000000111011    1011000000111100    1011000000111101    1011000000111110    1011000000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45115 - 45119

  --1011000001000000    1011000001000001    1011000001000010    1011000001000011    1011000001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45120 - 45124

  --1011000001000101    1011000001000110    1011000001000111    1011000001001000    1011000001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45125 - 45129

  --1011000001001010    1011000001001011    1011000001001100    1011000001001101    1011000001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45130 - 45134

  --1011000001001111    1011000001010000    1011000001010001    1011000001010010    1011000001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45135 - 45139

  --1011000001010100    1011000001010101    1011000001010110    1011000001010111    1011000001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45140 - 45144

  --1011000001011001    1011000001011010    1011000001011011    1011000001011100    1011000001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45145 - 45149

  --1011000001011110    1011000001011111    1011000001100000    1011000001100001    1011000001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45150 - 45154

  --1011000001100011    1011000001100100    1011000001100101    1011000001100110    1011000001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45155 - 45159

  --1011000001101000    1011000001101001    1011000001101010    1011000001101011    1011000001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45160 - 45164

  --1011000001101101    1011000001101110    1011000001101111    1011000001110000    1011000001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45165 - 45169

  --1011000001110010    1011000001110011    1011000001110100    1011000001110101    1011000001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45170 - 45174

  --1011000001110111    1011000001111000    1011000001111001    1011000001111010    1011000001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45175 - 45179

  --1011000001111100    1011000001111101    1011000001111110    1011000001111111    1011000010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45180 - 45184

  --1011000010000001    1011000010000010    1011000010000011    1011000010000100    1011000010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45185 - 45189

  --1011000010000110    1011000010000111    1011000010001000    1011000010001001    1011000010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45190 - 45194

  --1011000010001011    1011000010001100    1011000010001101    1011000010001110    1011000010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45195 - 45199

  --1011000010010000    1011000010010001    1011000010010010    1011000010010011    1011000010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45200 - 45204

  --1011000010010101    1011000010010110    1011000010010111    1011000010011000    1011000010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45205 - 45209

  --1011000010011010    1011000010011011    1011000010011100    1011000010011101    1011000010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45210 - 45214

  --1011000010011111    1011000010100000    1011000010100001    1011000010100010    1011000010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45215 - 45219

  --1011000010100100    1011000010100101    1011000010100110    1011000010100111    1011000010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45220 - 45224

  --1011000010101001    1011000010101010    1011000010101011    1011000010101100    1011000010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45225 - 45229

  --1011000010101110    1011000010101111    1011000010110000    1011000010110001    1011000010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45230 - 45234

  --1011000010110011    1011000010110100    1011000010110101    1011000010110110    1011000010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45235 - 45239

  --1011000010111000    1011000010111001    1011000010111010    1011000010111011    1011000010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45240 - 45244

  --1011000010111101    1011000010111110    1011000010111111    1011000011000000    1011000011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45245 - 45249

  --1011000011000010    1011000011000011    1011000011000100    1011000011000101    1011000011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45250 - 45254

  --1011000011000111    1011000011001000    1011000011001001    1011000011001010    1011000011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45255 - 45259

  --1011000011001100    1011000011001101    1011000011001110    1011000011001111    1011000011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45260 - 45264

  --1011000011010001    1011000011010010    1011000011010011    1011000011010100    1011000011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45265 - 45269

  --1011000011010110    1011000011010111    1011000011011000    1011000011011001    1011000011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45270 - 45274

  --1011000011011011    1011000011011100    1011000011011101    1011000011011110    1011000011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45275 - 45279

  --1011000011100000    1011000011100001    1011000011100010    1011000011100011    1011000011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45280 - 45284

  --1011000011100101    1011000011100110    1011000011100111    1011000011101000    1011000011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45285 - 45289

  --1011000011101010    1011000011101011    1011000011101100    1011000011101101    1011000011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45290 - 45294

  --1011000011101111    1011000011110000    1011000011110001    1011000011110010    1011000011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45295 - 45299

  --1011000011110100    1011000011110101    1011000011110110    1011000011110111    1011000011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45300 - 45304

  --1011000011111001    1011000011111010    1011000011111011    1011000011111100    1011000011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45305 - 45309

  --1011000011111110    1011000011111111    1011000100000000    1011000100000001    1011000100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45310 - 45314

  --1011000100000011    1011000100000100    1011000100000101    1011000100000110    1011000100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45315 - 45319

  --1011000100001000    1011000100001001    1011000100001010    1011000100001011    1011000100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45320 - 45324

  --1011000100001101    1011000100001110    1011000100001111    1011000100010000    1011000100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45325 - 45329

  --1011000100010010    1011000100010011    1011000100010100    1011000100010101    1011000100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45330 - 45334

  --1011000100010111    1011000100011000    1011000100011001    1011000100011010    1011000100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45335 - 45339

  --1011000100011100    1011000100011101    1011000100011110    1011000100011111    1011000100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45340 - 45344

  --1011000100100001    1011000100100010    1011000100100011    1011000100100100    1011000100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45345 - 45349

  --1011000100100110    1011000100100111    1011000100101000    1011000100101001    1011000100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45350 - 45354

  --1011000100101011    1011000100101100    1011000100101101    1011000100101110    1011000100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45355 - 45359

  --1011000100110000    1011000100110001    1011000100110010    1011000100110011    1011000100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45360 - 45364

  --1011000100110101    1011000100110110    1011000100110111    1011000100111000    1011000100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45365 - 45369

  --1011000100111010    1011000100111011    1011000100111100    1011000100111101    1011000100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45370 - 45374

  --1011000100111111    1011000101000000    1011000101000001    1011000101000010    1011000101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45375 - 45379

  --1011000101000100    1011000101000101    1011000101000110    1011000101000111    1011000101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45380 - 45384

  --1011000101001001    1011000101001010    1011000101001011    1011000101001100    1011000101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45385 - 45389

  --1011000101001110    1011000101001111    1011000101010000    1011000101010001    1011000101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45390 - 45394

  --1011000101010011    1011000101010100    1011000101010101    1011000101010110    1011000101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45395 - 45399

  --1011000101011000    1011000101011001    1011000101011010    1011000101011011    1011000101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45400 - 45404

  --1011000101011101    1011000101011110    1011000101011111    1011000101100000    1011000101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45405 - 45409

  --1011000101100010    1011000101100011    1011000101100100    1011000101100101    1011000101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45410 - 45414

  --1011000101100111    1011000101101000    1011000101101001    1011000101101010    1011000101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45415 - 45419

  --1011000101101100    1011000101101101    1011000101101110    1011000101101111    1011000101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45420 - 45424

  --1011000101110001    1011000101110010    1011000101110011    1011000101110100    1011000101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45425 - 45429

  --1011000101110110    1011000101110111    1011000101111000    1011000101111001    1011000101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45430 - 45434

  --1011000101111011    1011000101111100    1011000101111101    1011000101111110    1011000101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45435 - 45439

  --1011000110000000    1011000110000001    1011000110000010    1011000110000011    1011000110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45440 - 45444

  --1011000110000101    1011000110000110    1011000110000111    1011000110001000    1011000110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45445 - 45449

  --1011000110001010    1011000110001011    1011000110001100    1011000110001101    1011000110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45450 - 45454

  --1011000110001111    1011000110010000    1011000110010001    1011000110010010    1011000110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45455 - 45459

  --1011000110010100    1011000110010101    1011000110010110    1011000110010111    1011000110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45460 - 45464

  --1011000110011001    1011000110011010    1011000110011011    1011000110011100    1011000110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45465 - 45469

  --1011000110011110    1011000110011111    1011000110100000    1011000110100001    1011000110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45470 - 45474

  --1011000110100011    1011000110100100    1011000110100101    1011000110100110    1011000110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45475 - 45479

  --1011000110101000    1011000110101001    1011000110101010    1011000110101011    1011000110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45480 - 45484

  --1011000110101101    1011000110101110    1011000110101111    1011000110110000    1011000110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45485 - 45489

  --1011000110110010    1011000110110011    1011000110110100    1011000110110101    1011000110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45490 - 45494

  --1011000110110111    1011000110111000    1011000110111001    1011000110111010    1011000110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45495 - 45499

  --1011000110111100    1011000110111101    1011000110111110    1011000110111111    1011000111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45500 - 45504

  --1011000111000001    1011000111000010    1011000111000011    1011000111000100    1011000111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45505 - 45509

  --1011000111000110    1011000111000111    1011000111001000    1011000111001001    1011000111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45510 - 45514

  --1011000111001011    1011000111001100    1011000111001101    1011000111001110    1011000111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45515 - 45519

  --1011000111010000    1011000111010001    1011000111010010    1011000111010011    1011000111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45520 - 45524

  --1011000111010101    1011000111010110    1011000111010111    1011000111011000    1011000111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45525 - 45529

  --1011000111011010    1011000111011011    1011000111011100    1011000111011101    1011000111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45530 - 45534

  --1011000111011111    1011000111100000    1011000111100001    1011000111100010    1011000111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45535 - 45539

  --1011000111100100    1011000111100101    1011000111100110    1011000111100111    1011000111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45540 - 45544

  --1011000111101001    1011000111101010    1011000111101011    1011000111101100    1011000111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45545 - 45549

  --1011000111101110    1011000111101111    1011000111110000    1011000111110001    1011000111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45550 - 45554

  --1011000111110011    1011000111110100    1011000111110101    1011000111110110    1011000111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45555 - 45559

  --1011000111111000    1011000111111001    1011000111111010    1011000111111011    1011000111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45560 - 45564

  --1011000111111101    1011000111111110    1011000111111111    1011001000000000    1011001000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45565 - 45569

  --1011001000000010    1011001000000011    1011001000000100    1011001000000101    1011001000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45570 - 45574

  --1011001000000111    1011001000001000    1011001000001001    1011001000001010    1011001000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45575 - 45579

  --1011001000001100    1011001000001101    1011001000001110    1011001000001111    1011001000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45580 - 45584

  --1011001000010001    1011001000010010    1011001000010011    1011001000010100    1011001000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45585 - 45589

  --1011001000010110    1011001000010111    1011001000011000    1011001000011001    1011001000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45590 - 45594

  --1011001000011011    1011001000011100    1011001000011101    1011001000011110    1011001000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45595 - 45599

  --1011001000100000    1011001000100001    1011001000100010    1011001000100011    1011001000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45600 - 45604

  --1011001000100101    1011001000100110    1011001000100111    1011001000101000    1011001000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45605 - 45609

  --1011001000101010    1011001000101011    1011001000101100    1011001000101101    1011001000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45610 - 45614

  --1011001000101111    1011001000110000    1011001000110001    1011001000110010    1011001000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45615 - 45619

  --1011001000110100    1011001000110101    1011001000110110    1011001000110111    1011001000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45620 - 45624

  --1011001000111001    1011001000111010    1011001000111011    1011001000111100    1011001000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45625 - 45629

  --1011001000111110    1011001000111111    1011001001000000    1011001001000001    1011001001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45630 - 45634

  --1011001001000011    1011001001000100    1011001001000101    1011001001000110    1011001001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45635 - 45639

  --1011001001001000    1011001001001001    1011001001001010    1011001001001011    1011001001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45640 - 45644

  --1011001001001101    1011001001001110    1011001001001111    1011001001010000    1011001001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45645 - 45649

  --1011001001010010    1011001001010011    1011001001010100    1011001001010101    1011001001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45650 - 45654

  --1011001001010111    1011001001011000    1011001001011001    1011001001011010    1011001001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45655 - 45659

  --1011001001011100    1011001001011101    1011001001011110    1011001001011111    1011001001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45660 - 45664

  --1011001001100001    1011001001100010    1011001001100011    1011001001100100    1011001001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45665 - 45669

  --1011001001100110    1011001001100111    1011001001101000    1011001001101001    1011001001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45670 - 45674

  --1011001001101011    1011001001101100    1011001001101101    1011001001101110    1011001001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45675 - 45679

  --1011001001110000    1011001001110001    1011001001110010    1011001001110011    1011001001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45680 - 45684

  --1011001001110101    1011001001110110    1011001001110111    1011001001111000    1011001001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45685 - 45689

  --1011001001111010    1011001001111011    1011001001111100    1011001001111101    1011001001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45690 - 45694

  --1011001001111111    1011001010000000    1011001010000001    1011001010000010    1011001010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45695 - 45699

  --1011001010000100    1011001010000101    1011001010000110    1011001010000111    1011001010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45700 - 45704

  --1011001010001001    1011001010001010    1011001010001011    1011001010001100    1011001010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45705 - 45709

  --1011001010001110    1011001010001111    1011001010010000    1011001010010001    1011001010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45710 - 45714

  --1011001010010011    1011001010010100    1011001010010101    1011001010010110    1011001010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45715 - 45719

  --1011001010011000    1011001010011001    1011001010011010    1011001010011011    1011001010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45720 - 45724

  --1011001010011101    1011001010011110    1011001010011111    1011001010100000    1011001010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45725 - 45729

  --1011001010100010    1011001010100011    1011001010100100    1011001010100101    1011001010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45730 - 45734

  --1011001010100111    1011001010101000    1011001010101001    1011001010101010    1011001010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45735 - 45739

  --1011001010101100    1011001010101101    1011001010101110    1011001010101111    1011001010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45740 - 45744

  --1011001010110001    1011001010110010    1011001010110011    1011001010110100    1011001010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45745 - 45749

  --1011001010110110    1011001010110111    1011001010111000    1011001010111001    1011001010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45750 - 45754

  --1011001010111011    1011001010111100    1011001010111101    1011001010111110    1011001010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45755 - 45759

  --1011001011000000    1011001011000001    1011001011000010    1011001011000011    1011001011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45760 - 45764

  --1011001011000101    1011001011000110    1011001011000111    1011001011001000    1011001011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45765 - 45769

  --1011001011001010    1011001011001011    1011001011001100    1011001011001101    1011001011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45770 - 45774

  --1011001011001111    1011001011010000    1011001011010001    1011001011010010    1011001011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45775 - 45779

  --1011001011010100    1011001011010101    1011001011010110    1011001011010111    1011001011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45780 - 45784

  --1011001011011001    1011001011011010    1011001011011011    1011001011011100    1011001011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45785 - 45789

  --1011001011011110    1011001011011111    1011001011100000    1011001011100001    1011001011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45790 - 45794

  --1011001011100011    1011001011100100    1011001011100101    1011001011100110    1011001011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45795 - 45799

  --1011001011101000    1011001011101001    1011001011101010    1011001011101011    1011001011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45800 - 45804

  --1011001011101101    1011001011101110    1011001011101111    1011001011110000    1011001011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45805 - 45809

  --1011001011110010    1011001011110011    1011001011110100    1011001011110101    1011001011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45810 - 45814

  --1011001011110111    1011001011111000    1011001011111001    1011001011111010    1011001011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45815 - 45819

  --1011001011111100    1011001011111101    1011001011111110    1011001011111111    1011001100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45820 - 45824

  --1011001100000001    1011001100000010    1011001100000011    1011001100000100    1011001100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45825 - 45829

  --1011001100000110    1011001100000111    1011001100001000    1011001100001001    1011001100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45830 - 45834

  --1011001100001011    1011001100001100    1011001100001101    1011001100001110    1011001100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45835 - 45839

  --1011001100010000    1011001100010001    1011001100010010    1011001100010011    1011001100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45840 - 45844

  --1011001100010101    1011001100010110    1011001100010111    1011001100011000    1011001100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45845 - 45849

  --1011001100011010    1011001100011011    1011001100011100    1011001100011101    1011001100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45850 - 45854

  --1011001100011111    1011001100100000    1011001100100001    1011001100100010    1011001100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45855 - 45859

  --1011001100100100    1011001100100101    1011001100100110    1011001100100111    1011001100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45860 - 45864

  --1011001100101001    1011001100101010    1011001100101011    1011001100101100    1011001100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45865 - 45869

  --1011001100101110    1011001100101111    1011001100110000    1011001100110001    1011001100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45870 - 45874

  --1011001100110011    1011001100110100    1011001100110101    1011001100110110    1011001100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45875 - 45879

  --1011001100111000    1011001100111001    1011001100111010    1011001100111011    1011001100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45880 - 45884

  --1011001100111101    1011001100111110    1011001100111111    1011001101000000    1011001101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45885 - 45889

  --1011001101000010    1011001101000011    1011001101000100    1011001101000101    1011001101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45890 - 45894

  --1011001101000111    1011001101001000    1011001101001001    1011001101001010    1011001101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45895 - 45899

  --1011001101001100    1011001101001101    1011001101001110    1011001101001111    1011001101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45900 - 45904

  --1011001101010001    1011001101010010    1011001101010011    1011001101010100    1011001101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45905 - 45909

  --1011001101010110    1011001101010111    1011001101011000    1011001101011001    1011001101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45910 - 45914

  --1011001101011011    1011001101011100    1011001101011101    1011001101011110    1011001101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45915 - 45919

  --1011001101100000    1011001101100001    1011001101100010    1011001101100011    1011001101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45920 - 45924

  --1011001101100101    1011001101100110    1011001101100111    1011001101101000    1011001101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45925 - 45929

  --1011001101101010    1011001101101011    1011001101101100    1011001101101101    1011001101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45930 - 45934

  --1011001101101111    1011001101110000    1011001101110001    1011001101110010    1011001101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45935 - 45939

  --1011001101110100    1011001101110101    1011001101110110    1011001101110111    1011001101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45940 - 45944

  --1011001101111001    1011001101111010    1011001101111011    1011001101111100    1011001101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45945 - 45949

  --1011001101111110    1011001101111111    1011001110000000    1011001110000001    1011001110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45950 - 45954

  --1011001110000011    1011001110000100    1011001110000101    1011001110000110    1011001110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45955 - 45959

  --1011001110001000    1011001110001001    1011001110001010    1011001110001011    1011001110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45960 - 45964

  --1011001110001101    1011001110001110    1011001110001111    1011001110010000    1011001110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45965 - 45969

  --1011001110010010    1011001110010011    1011001110010100    1011001110010101    1011001110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45970 - 45974

  --1011001110010111    1011001110011000    1011001110011001    1011001110011010    1011001110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45975 - 45979

  --1011001110011100    1011001110011101    1011001110011110    1011001110011111    1011001110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45980 - 45984

  --1011001110100001    1011001110100010    1011001110100011    1011001110100100    1011001110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45985 - 45989

  --1011001110100110    1011001110100111    1011001110101000    1011001110101001    1011001110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45990 - 45994

  --1011001110101011    1011001110101100    1011001110101101    1011001110101110    1011001110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 45995 - 45999

  --1011001110110000    1011001110110001    1011001110110010    1011001110110011    1011001110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46000 - 46004

  --1011001110110101    1011001110110110    1011001110110111    1011001110111000    1011001110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46005 - 46009

  --1011001110111010    1011001110111011    1011001110111100    1011001110111101    1011001110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46010 - 46014

  --1011001110111111    1011001111000000    1011001111000001    1011001111000010    1011001111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46015 - 46019

  --1011001111000100    1011001111000101    1011001111000110    1011001111000111    1011001111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46020 - 46024

  --1011001111001001    1011001111001010    1011001111001011    1011001111001100    1011001111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46025 - 46029

  --1011001111001110    1011001111001111    1011001111010000    1011001111010001    1011001111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46030 - 46034

  --1011001111010011    1011001111010100    1011001111010101    1011001111010110    1011001111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46035 - 46039

  --1011001111011000    1011001111011001    1011001111011010    1011001111011011    1011001111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46040 - 46044

  --1011001111011101    1011001111011110    1011001111011111    1011001111100000    1011001111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46045 - 46049

  --1011001111100010    1011001111100011    1011001111100100    1011001111100101    1011001111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46050 - 46054

  --1011001111100111    1011001111101000    1011001111101001    1011001111101010    1011001111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46055 - 46059

  --1011001111101100    1011001111101101    1011001111101110    1011001111101111    1011001111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46060 - 46064

  --1011001111110001    1011001111110010    1011001111110011    1011001111110100    1011001111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46065 - 46069

  --1011001111110110    1011001111110111    1011001111111000    1011001111111001    1011001111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46070 - 46074

  --1011001111111011    1011001111111100    1011001111111101    1011001111111110    1011001111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46075 - 46079

  --1011010000000000    1011010000000001    1011010000000010    1011010000000011    1011010000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46080 - 46084

  --1011010000000101    1011010000000110    1011010000000111    1011010000001000    1011010000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46085 - 46089

  --1011010000001010    1011010000001011    1011010000001100    1011010000001101    1011010000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46090 - 46094

  --1011010000001111    1011010000010000    1011010000010001    1011010000010010    1011010000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46095 - 46099

  --1011010000010100    1011010000010101    1011010000010110    1011010000010111    1011010000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46100 - 46104

  --1011010000011001    1011010000011010    1011010000011011    1011010000011100    1011010000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46105 - 46109

  --1011010000011110    1011010000011111    1011010000100000    1011010000100001    1011010000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46110 - 46114

  --1011010000100011    1011010000100100    1011010000100101    1011010000100110    1011010000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46115 - 46119

  --1011010000101000    1011010000101001    1011010000101010    1011010000101011    1011010000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46120 - 46124

  --1011010000101101    1011010000101110    1011010000101111    1011010000110000    1011010000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46125 - 46129

  --1011010000110010    1011010000110011    1011010000110100    1011010000110101    1011010000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46130 - 46134

  --1011010000110111    1011010000111000    1011010000111001    1011010000111010    1011010000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46135 - 46139

  --1011010000111100    1011010000111101    1011010000111110    1011010000111111    1011010001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46140 - 46144

  --1011010001000001    1011010001000010    1011010001000011    1011010001000100    1011010001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46145 - 46149

  --1011010001000110    1011010001000111    1011010001001000    1011010001001001    1011010001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46150 - 46154

  --1011010001001011    1011010001001100    1011010001001101    1011010001001110    1011010001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46155 - 46159

  --1011010001010000    1011010001010001    1011010001010010    1011010001010011    1011010001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46160 - 46164

  --1011010001010101    1011010001010110    1011010001010111    1011010001011000    1011010001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46165 - 46169

  --1011010001011010    1011010001011011    1011010001011100    1011010001011101    1011010001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46170 - 46174

  --1011010001011111    1011010001100000    1011010001100001    1011010001100010    1011010001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46175 - 46179

  --1011010001100100    1011010001100101    1011010001100110    1011010001100111    1011010001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46180 - 46184

  --1011010001101001    1011010001101010    1011010001101011    1011010001101100    1011010001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46185 - 46189

  --1011010001101110    1011010001101111    1011010001110000    1011010001110001    1011010001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46190 - 46194

  --1011010001110011    1011010001110100    1011010001110101    1011010001110110    1011010001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46195 - 46199

  --1011010001111000    1011010001111001    1011010001111010    1011010001111011    1011010001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46200 - 46204

  --1011010001111101    1011010001111110    1011010001111111    1011010010000000    1011010010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46205 - 46209

  --1011010010000010    1011010010000011    1011010010000100    1011010010000101    1011010010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46210 - 46214

  --1011010010000111    1011010010001000    1011010010001001    1011010010001010    1011010010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46215 - 46219

  --1011010010001100    1011010010001101    1011010010001110    1011010010001111    1011010010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46220 - 46224

  --1011010010010001    1011010010010010    1011010010010011    1011010010010100    1011010010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46225 - 46229

  --1011010010010110    1011010010010111    1011010010011000    1011010010011001    1011010010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46230 - 46234

  --1011010010011011    1011010010011100    1011010010011101    1011010010011110    1011010010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46235 - 46239

  --1011010010100000    1011010010100001    1011010010100010    1011010010100011    1011010010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46240 - 46244

  --1011010010100101    1011010010100110    1011010010100111    1011010010101000    1011010010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46245 - 46249

  --1011010010101010    1011010010101011    1011010010101100    1011010010101101    1011010010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46250 - 46254

  --1011010010101111    1011010010110000    1011010010110001    1011010010110010    1011010010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46255 - 46259

  --1011010010110100    1011010010110101    1011010010110110    1011010010110111    1011010010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46260 - 46264

  --1011010010111001    1011010010111010    1011010010111011    1011010010111100    1011010010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46265 - 46269

  --1011010010111110    1011010010111111    1011010011000000    1011010011000001    1011010011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46270 - 46274

  --1011010011000011    1011010011000100    1011010011000101    1011010011000110    1011010011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46275 - 46279

  --1011010011001000    1011010011001001    1011010011001010    1011010011001011    1011010011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46280 - 46284

  --1011010011001101    1011010011001110    1011010011001111    1011010011010000    1011010011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46285 - 46289

  --1011010011010010    1011010011010011    1011010011010100    1011010011010101    1011010011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46290 - 46294

  --1011010011010111    1011010011011000    1011010011011001    1011010011011010    1011010011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46295 - 46299

  --1011010011011100    1011010011011101    1011010011011110    1011010011011111    1011010011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46300 - 46304

  --1011010011100001    1011010011100010    1011010011100011    1011010011100100    1011010011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46305 - 46309

  --1011010011100110    1011010011100111    1011010011101000    1011010011101001    1011010011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46310 - 46314

  --1011010011101011    1011010011101100    1011010011101101    1011010011101110    1011010011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46315 - 46319

  --1011010011110000    1011010011110001    1011010011110010    1011010011110011    1011010011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46320 - 46324

  --1011010011110101    1011010011110110    1011010011110111    1011010011111000    1011010011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46325 - 46329

  --1011010011111010    1011010011111011    1011010011111100    1011010011111101    1011010011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46330 - 46334

  --1011010011111111    1011010100000000    1011010100000001    1011010100000010    1011010100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46335 - 46339

  --1011010100000100    1011010100000101    1011010100000110    1011010100000111    1011010100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46340 - 46344

  --1011010100001001    1011010100001010    1011010100001011    1011010100001100    1011010100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46345 - 46349

  --1011010100001110    1011010100001111    1011010100010000    1011010100010001    1011010100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46350 - 46354

  --1011010100010011    1011010100010100    1011010100010101    1011010100010110    1011010100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46355 - 46359

  --1011010100011000    1011010100011001    1011010100011010    1011010100011011    1011010100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46360 - 46364

  --1011010100011101    1011010100011110    1011010100011111    1011010100100000    1011010100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46365 - 46369

  --1011010100100010    1011010100100011    1011010100100100    1011010100100101    1011010100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46370 - 46374

  --1011010100100111    1011010100101000    1011010100101001    1011010100101010    1011010100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46375 - 46379

  --1011010100101100    1011010100101101    1011010100101110    1011010100101111    1011010100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46380 - 46384

  --1011010100110001    1011010100110010    1011010100110011    1011010100110100    1011010100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46385 - 46389

  --1011010100110110    1011010100110111    1011010100111000    1011010100111001    1011010100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46390 - 46394

  --1011010100111011    1011010100111100    1011010100111101    1011010100111110    1011010100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46395 - 46399

  --1011010101000000    1011010101000001    1011010101000010    1011010101000011    1011010101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46400 - 46404

  --1011010101000101    1011010101000110    1011010101000111    1011010101001000    1011010101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46405 - 46409

  --1011010101001010    1011010101001011    1011010101001100    1011010101001101    1011010101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46410 - 46414

  --1011010101001111    1011010101010000    1011010101010001    1011010101010010    1011010101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46415 - 46419

  --1011010101010100    1011010101010101    1011010101010110    1011010101010111    1011010101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46420 - 46424

  --1011010101011001    1011010101011010    1011010101011011    1011010101011100    1011010101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46425 - 46429

  --1011010101011110    1011010101011111    1011010101100000    1011010101100001    1011010101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46430 - 46434

  --1011010101100011    1011010101100100    1011010101100101    1011010101100110    1011010101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46435 - 46439

  --1011010101101000    1011010101101001    1011010101101010    1011010101101011    1011010101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46440 - 46444

  --1011010101101101    1011010101101110    1011010101101111    1011010101110000    1011010101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46445 - 46449

  --1011010101110010    1011010101110011    1011010101110100    1011010101110101    1011010101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46450 - 46454

  --1011010101110111    1011010101111000    1011010101111001    1011010101111010    1011010101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46455 - 46459

  --1011010101111100    1011010101111101    1011010101111110    1011010101111111    1011010110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46460 - 46464

  --1011010110000001    1011010110000010    1011010110000011    1011010110000100    1011010110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46465 - 46469

  --1011010110000110    1011010110000111    1011010110001000    1011010110001001    1011010110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46470 - 46474

  --1011010110001011    1011010110001100    1011010110001101    1011010110001110    1011010110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46475 - 46479

  --1011010110010000    1011010110010001    1011010110010010    1011010110010011    1011010110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46480 - 46484

  --1011010110010101    1011010110010110    1011010110010111    1011010110011000    1011010110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46485 - 46489

  --1011010110011010    1011010110011011    1011010110011100    1011010110011101    1011010110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46490 - 46494

  --1011010110011111    1011010110100000    1011010110100001    1011010110100010    1011010110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46495 - 46499

  --1011010110100100    1011010110100101    1011010110100110    1011010110100111    1011010110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46500 - 46504

  --1011010110101001    1011010110101010    1011010110101011    1011010110101100    1011010110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46505 - 46509

  --1011010110101110    1011010110101111    1011010110110000    1011010110110001    1011010110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46510 - 46514

  --1011010110110011    1011010110110100    1011010110110101    1011010110110110    1011010110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46515 - 46519

  --1011010110111000    1011010110111001    1011010110111010    1011010110111011    1011010110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46520 - 46524

  --1011010110111101    1011010110111110    1011010110111111    1011010111000000    1011010111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46525 - 46529

  --1011010111000010    1011010111000011    1011010111000100    1011010111000101    1011010111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46530 - 46534

  --1011010111000111    1011010111001000    1011010111001001    1011010111001010    1011010111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46535 - 46539

  --1011010111001100    1011010111001101    1011010111001110    1011010111001111    1011010111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46540 - 46544

  --1011010111010001    1011010111010010    1011010111010011    1011010111010100    1011010111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46545 - 46549

  --1011010111010110    1011010111010111    1011010111011000    1011010111011001    1011010111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46550 - 46554

  --1011010111011011    1011010111011100    1011010111011101    1011010111011110    1011010111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46555 - 46559

  --1011010111100000    1011010111100001    1011010111100010    1011010111100011    1011010111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46560 - 46564

  --1011010111100101    1011010111100110    1011010111100111    1011010111101000    1011010111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46565 - 46569

  --1011010111101010    1011010111101011    1011010111101100    1011010111101101    1011010111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46570 - 46574

  --1011010111101111    1011010111110000    1011010111110001    1011010111110010    1011010111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46575 - 46579

  --1011010111110100    1011010111110101    1011010111110110    1011010111110111    1011010111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46580 - 46584

  --1011010111111001    1011010111111010    1011010111111011    1011010111111100    1011010111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46585 - 46589

  --1011010111111110    1011010111111111    1011011000000000    1011011000000001    1011011000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46590 - 46594

  --1011011000000011    1011011000000100    1011011000000101    1011011000000110    1011011000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46595 - 46599

  --1011011000001000    1011011000001001    1011011000001010    1011011000001011    1011011000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46600 - 46604

  --1011011000001101    1011011000001110    1011011000001111    1011011000010000    1011011000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46605 - 46609

  --1011011000010010    1011011000010011    1011011000010100    1011011000010101    1011011000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46610 - 46614

  --1011011000010111    1011011000011000    1011011000011001    1011011000011010    1011011000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46615 - 46619

  --1011011000011100    1011011000011101    1011011000011110    1011011000011111    1011011000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46620 - 46624

  --1011011000100001    1011011000100010    1011011000100011    1011011000100100    1011011000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46625 - 46629

  --1011011000100110    1011011000100111    1011011000101000    1011011000101001    1011011000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46630 - 46634

  --1011011000101011    1011011000101100    1011011000101101    1011011000101110    1011011000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46635 - 46639

  --1011011000110000    1011011000110001    1011011000110010    1011011000110011    1011011000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46640 - 46644

  --1011011000110101    1011011000110110    1011011000110111    1011011000111000    1011011000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46645 - 46649

  --1011011000111010    1011011000111011    1011011000111100    1011011000111101    1011011000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46650 - 46654

  --1011011000111111    1011011001000000    1011011001000001    1011011001000010    1011011001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46655 - 46659

  --1011011001000100    1011011001000101    1011011001000110    1011011001000111    1011011001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46660 - 46664

  --1011011001001001    1011011001001010    1011011001001011    1011011001001100    1011011001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46665 - 46669

  --1011011001001110    1011011001001111    1011011001010000    1011011001010001    1011011001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46670 - 46674

  --1011011001010011    1011011001010100    1011011001010101    1011011001010110    1011011001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46675 - 46679

  --1011011001011000    1011011001011001    1011011001011010    1011011001011011    1011011001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46680 - 46684

  --1011011001011101    1011011001011110    1011011001011111    1011011001100000    1011011001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46685 - 46689

  --1011011001100010    1011011001100011    1011011001100100    1011011001100101    1011011001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46690 - 46694

  --1011011001100111    1011011001101000    1011011001101001    1011011001101010    1011011001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46695 - 46699

  --1011011001101100    1011011001101101    1011011001101110    1011011001101111    1011011001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46700 - 46704

  --1011011001110001    1011011001110010    1011011001110011    1011011001110100    1011011001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46705 - 46709

  --1011011001110110    1011011001110111    1011011001111000    1011011001111001    1011011001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46710 - 46714

  --1011011001111011    1011011001111100    1011011001111101    1011011001111110    1011011001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46715 - 46719

  --1011011010000000    1011011010000001    1011011010000010    1011011010000011    1011011010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46720 - 46724

  --1011011010000101    1011011010000110    1011011010000111    1011011010001000    1011011010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46725 - 46729

  --1011011010001010    1011011010001011    1011011010001100    1011011010001101    1011011010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46730 - 46734

  --1011011010001111    1011011010010000    1011011010010001    1011011010010010    1011011010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46735 - 46739

  --1011011010010100    1011011010010101    1011011010010110    1011011010010111    1011011010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46740 - 46744

  --1011011010011001    1011011010011010    1011011010011011    1011011010011100    1011011010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46745 - 46749

  --1011011010011110    1011011010011111    1011011010100000    1011011010100001    1011011010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46750 - 46754

  --1011011010100011    1011011010100100    1011011010100101    1011011010100110    1011011010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46755 - 46759

  --1011011010101000    1011011010101001    1011011010101010    1011011010101011    1011011010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46760 - 46764

  --1011011010101101    1011011010101110    1011011010101111    1011011010110000    1011011010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46765 - 46769

  --1011011010110010    1011011010110011    1011011010110100    1011011010110101    1011011010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46770 - 46774

  --1011011010110111    1011011010111000    1011011010111001    1011011010111010    1011011010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46775 - 46779

  --1011011010111100    1011011010111101    1011011010111110    1011011010111111    1011011011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46780 - 46784

  --1011011011000001    1011011011000010    1011011011000011    1011011011000100    1011011011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46785 - 46789

  --1011011011000110    1011011011000111    1011011011001000    1011011011001001    1011011011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46790 - 46794

  --1011011011001011    1011011011001100    1011011011001101    1011011011001110    1011011011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46795 - 46799

  --1011011011010000    1011011011010001    1011011011010010    1011011011010011    1011011011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46800 - 46804

  --1011011011010101    1011011011010110    1011011011010111    1011011011011000    1011011011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46805 - 46809

  --1011011011011010    1011011011011011    1011011011011100    1011011011011101    1011011011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46810 - 46814

  --1011011011011111    1011011011100000    1011011011100001    1011011011100010    1011011011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46815 - 46819

  --1011011011100100    1011011011100101    1011011011100110    1011011011100111    1011011011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46820 - 46824

  --1011011011101001    1011011011101010    1011011011101011    1011011011101100    1011011011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46825 - 46829

  --1011011011101110    1011011011101111    1011011011110000    1011011011110001    1011011011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46830 - 46834

  --1011011011110011    1011011011110100    1011011011110101    1011011011110110    1011011011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46835 - 46839

  --1011011011111000    1011011011111001    1011011011111010    1011011011111011    1011011011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46840 - 46844

  --1011011011111101    1011011011111110    1011011011111111    1011011100000000    1011011100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46845 - 46849

  --1011011100000010    1011011100000011    1011011100000100    1011011100000101    1011011100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46850 - 46854

  --1011011100000111    1011011100001000    1011011100001001    1011011100001010    1011011100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46855 - 46859

  --1011011100001100    1011011100001101    1011011100001110    1011011100001111    1011011100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46860 - 46864

  --1011011100010001    1011011100010010    1011011100010011    1011011100010100    1011011100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46865 - 46869

  --1011011100010110    1011011100010111    1011011100011000    1011011100011001    1011011100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46870 - 46874

  --1011011100011011    1011011100011100    1011011100011101    1011011100011110    1011011100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46875 - 46879

  --1011011100100000    1011011100100001    1011011100100010    1011011100100011    1011011100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46880 - 46884

  --1011011100100101    1011011100100110    1011011100100111    1011011100101000    1011011100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46885 - 46889

  --1011011100101010    1011011100101011    1011011100101100    1011011100101101    1011011100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46890 - 46894

  --1011011100101111    1011011100110000    1011011100110001    1011011100110010    1011011100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46895 - 46899

  --1011011100110100    1011011100110101    1011011100110110    1011011100110111    1011011100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46900 - 46904

  --1011011100111001    1011011100111010    1011011100111011    1011011100111100    1011011100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46905 - 46909

  --1011011100111110    1011011100111111    1011011101000000    1011011101000001    1011011101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46910 - 46914

  --1011011101000011    1011011101000100    1011011101000101    1011011101000110    1011011101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46915 - 46919

  --1011011101001000    1011011101001001    1011011101001010    1011011101001011    1011011101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46920 - 46924

  --1011011101001101    1011011101001110    1011011101001111    1011011101010000    1011011101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46925 - 46929

  --1011011101010010    1011011101010011    1011011101010100    1011011101010101    1011011101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46930 - 46934

  --1011011101010111    1011011101011000    1011011101011001    1011011101011010    1011011101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46935 - 46939

  --1011011101011100    1011011101011101    1011011101011110    1011011101011111    1011011101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46940 - 46944

  --1011011101100001    1011011101100010    1011011101100011    1011011101100100    1011011101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46945 - 46949

  --1011011101100110    1011011101100111    1011011101101000    1011011101101001    1011011101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46950 - 46954

  --1011011101101011    1011011101101100    1011011101101101    1011011101101110    1011011101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46955 - 46959

  --1011011101110000    1011011101110001    1011011101110010    1011011101110011    1011011101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46960 - 46964

  --1011011101110101    1011011101110110    1011011101110111    1011011101111000    1011011101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46965 - 46969

  --1011011101111010    1011011101111011    1011011101111100    1011011101111101    1011011101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46970 - 46974

  --1011011101111111    1011011110000000    1011011110000001    1011011110000010    1011011110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46975 - 46979

  --1011011110000100    1011011110000101    1011011110000110    1011011110000111    1011011110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46980 - 46984

  --1011011110001001    1011011110001010    1011011110001011    1011011110001100    1011011110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46985 - 46989

  --1011011110001110    1011011110001111    1011011110010000    1011011110010001    1011011110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46990 - 46994

  --1011011110010011    1011011110010100    1011011110010101    1011011110010110    1011011110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 46995 - 46999

  --1011011110011000    1011011110011001    1011011110011010    1011011110011011    1011011110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47000 - 47004

  --1011011110011101    1011011110011110    1011011110011111    1011011110100000    1011011110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47005 - 47009

  --1011011110100010    1011011110100011    1011011110100100    1011011110100101    1011011110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47010 - 47014

  --1011011110100111    1011011110101000    1011011110101001    1011011110101010    1011011110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47015 - 47019

  --1011011110101100    1011011110101101    1011011110101110    1011011110101111    1011011110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47020 - 47024

  --1011011110110001    1011011110110010    1011011110110011    1011011110110100    1011011110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47025 - 47029

  --1011011110110110    1011011110110111    1011011110111000    1011011110111001    1011011110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47030 - 47034

  --1011011110111011    1011011110111100    1011011110111101    1011011110111110    1011011110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47035 - 47039

  --1011011111000000    1011011111000001    1011011111000010    1011011111000011    1011011111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47040 - 47044

  --1011011111000101    1011011111000110    1011011111000111    1011011111001000    1011011111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47045 - 47049

  --1011011111001010    1011011111001011    1011011111001100    1011011111001101    1011011111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47050 - 47054

  --1011011111001111    1011011111010000    1011011111010001    1011011111010010    1011011111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47055 - 47059

  --1011011111010100    1011011111010101    1011011111010110    1011011111010111    1011011111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47060 - 47064

  --1011011111011001    1011011111011010    1011011111011011    1011011111011100    1011011111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47065 - 47069

  --1011011111011110    1011011111011111    1011011111100000    1011011111100001    1011011111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47070 - 47074

  --1011011111100011    1011011111100100    1011011111100101    1011011111100110    1011011111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47075 - 47079

  --1011011111101000    1011011111101001    1011011111101010    1011011111101011    1011011111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47080 - 47084

  --1011011111101101    1011011111101110    1011011111101111    1011011111110000    1011011111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47085 - 47089

  --1011011111110010    1011011111110011    1011011111110100    1011011111110101    1011011111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47090 - 47094

  --1011011111110111    1011011111111000    1011011111111001    1011011111111010    1011011111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47095 - 47099

  --1011011111111100    1011011111111101    1011011111111110    1011011111111111    1011100000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47100 - 47104

  --1011100000000001    1011100000000010    1011100000000011    1011100000000100    1011100000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47105 - 47109

  --1011100000000110    1011100000000111    1011100000001000    1011100000001001    1011100000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47110 - 47114

  --1011100000001011    1011100000001100    1011100000001101    1011100000001110    1011100000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47115 - 47119

  --1011100000010000    1011100000010001    1011100000010010    1011100000010011    1011100000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47120 - 47124

  --1011100000010101    1011100000010110    1011100000010111    1011100000011000    1011100000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47125 - 47129

  --1011100000011010    1011100000011011    1011100000011100    1011100000011101    1011100000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47130 - 47134

  --1011100000011111    1011100000100000    1011100000100001    1011100000100010    1011100000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47135 - 47139

  --1011100000100100    1011100000100101    1011100000100110    1011100000100111    1011100000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47140 - 47144

  --1011100000101001    1011100000101010    1011100000101011    1011100000101100    1011100000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47145 - 47149

  --1011100000101110    1011100000101111    1011100000110000    1011100000110001    1011100000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47150 - 47154

  --1011100000110011    1011100000110100    1011100000110101    1011100000110110    1011100000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47155 - 47159

  --1011100000111000    1011100000111001    1011100000111010    1011100000111011    1011100000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47160 - 47164

  --1011100000111101    1011100000111110    1011100000111111    1011100001000000    1011100001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47165 - 47169

  --1011100001000010    1011100001000011    1011100001000100    1011100001000101    1011100001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47170 - 47174

  --1011100001000111    1011100001001000    1011100001001001    1011100001001010    1011100001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47175 - 47179

  --1011100001001100    1011100001001101    1011100001001110    1011100001001111    1011100001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47180 - 47184

  --1011100001010001    1011100001010010    1011100001010011    1011100001010100    1011100001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47185 - 47189

  --1011100001010110    1011100001010111    1011100001011000    1011100001011001    1011100001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47190 - 47194

  --1011100001011011    1011100001011100    1011100001011101    1011100001011110    1011100001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47195 - 47199

  --1011100001100000    1011100001100001    1011100001100010    1011100001100011    1011100001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47200 - 47204

  --1011100001100101    1011100001100110    1011100001100111    1011100001101000    1011100001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47205 - 47209

  --1011100001101010    1011100001101011    1011100001101100    1011100001101101    1011100001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47210 - 47214

  --1011100001101111    1011100001110000    1011100001110001    1011100001110010    1011100001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47215 - 47219

  --1011100001110100    1011100001110101    1011100001110110    1011100001110111    1011100001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47220 - 47224

  --1011100001111001    1011100001111010    1011100001111011    1011100001111100    1011100001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47225 - 47229

  --1011100001111110    1011100001111111    1011100010000000    1011100010000001    1011100010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47230 - 47234

  --1011100010000011    1011100010000100    1011100010000101    1011100010000110    1011100010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47235 - 47239

  --1011100010001000    1011100010001001    1011100010001010    1011100010001011    1011100010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47240 - 47244

  --1011100010001101    1011100010001110    1011100010001111    1011100010010000    1011100010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47245 - 47249

  --1011100010010010    1011100010010011    1011100010010100    1011100010010101    1011100010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47250 - 47254

  --1011100010010111    1011100010011000    1011100010011001    1011100010011010    1011100010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47255 - 47259

  --1011100010011100    1011100010011101    1011100010011110    1011100010011111    1011100010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47260 - 47264

  --1011100010100001    1011100010100010    1011100010100011    1011100010100100    1011100010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47265 - 47269

  --1011100010100110    1011100010100111    1011100010101000    1011100010101001    1011100010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47270 - 47274

  --1011100010101011    1011100010101100    1011100010101101    1011100010101110    1011100010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47275 - 47279

  --1011100010110000    1011100010110001    1011100010110010    1011100010110011    1011100010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47280 - 47284

  --1011100010110101    1011100010110110    1011100010110111    1011100010111000    1011100010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47285 - 47289

  --1011100010111010    1011100010111011    1011100010111100    1011100010111101    1011100010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47290 - 47294

  --1011100010111111    1011100011000000    1011100011000001    1011100011000010    1011100011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47295 - 47299

  --1011100011000100    1011100011000101    1011100011000110    1011100011000111    1011100011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47300 - 47304

  --1011100011001001    1011100011001010    1011100011001011    1011100011001100    1011100011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47305 - 47309

  --1011100011001110    1011100011001111    1011100011010000    1011100011010001    1011100011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47310 - 47314

  --1011100011010011    1011100011010100    1011100011010101    1011100011010110    1011100011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47315 - 47319

  --1011100011011000    1011100011011001    1011100011011010    1011100011011011    1011100011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47320 - 47324

  --1011100011011101    1011100011011110    1011100011011111    1011100011100000    1011100011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47325 - 47329

  --1011100011100010    1011100011100011    1011100011100100    1011100011100101    1011100011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47330 - 47334

  --1011100011100111    1011100011101000    1011100011101001    1011100011101010    1011100011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47335 - 47339

  --1011100011101100    1011100011101101    1011100011101110    1011100011101111    1011100011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47340 - 47344

  --1011100011110001    1011100011110010    1011100011110011    1011100011110100    1011100011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47345 - 47349

  --1011100011110110    1011100011110111    1011100011111000    1011100011111001    1011100011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47350 - 47354

  --1011100011111011    1011100011111100    1011100011111101    1011100011111110    1011100011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47355 - 47359

  --1011100100000000    1011100100000001    1011100100000010    1011100100000011    1011100100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47360 - 47364

  --1011100100000101    1011100100000110    1011100100000111    1011100100001000    1011100100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47365 - 47369

  --1011100100001010    1011100100001011    1011100100001100    1011100100001101    1011100100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47370 - 47374

  --1011100100001111    1011100100010000    1011100100010001    1011100100010010    1011100100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47375 - 47379

  --1011100100010100    1011100100010101    1011100100010110    1011100100010111    1011100100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47380 - 47384

  --1011100100011001    1011100100011010    1011100100011011    1011100100011100    1011100100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47385 - 47389

  --1011100100011110    1011100100011111    1011100100100000    1011100100100001    1011100100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47390 - 47394

  --1011100100100011    1011100100100100    1011100100100101    1011100100100110    1011100100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47395 - 47399

  --1011100100101000    1011100100101001    1011100100101010    1011100100101011    1011100100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47400 - 47404

  --1011100100101101    1011100100101110    1011100100101111    1011100100110000    1011100100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47405 - 47409

  --1011100100110010    1011100100110011    1011100100110100    1011100100110101    1011100100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47410 - 47414

  --1011100100110111    1011100100111000    1011100100111001    1011100100111010    1011100100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47415 - 47419

  --1011100100111100    1011100100111101    1011100100111110    1011100100111111    1011100101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47420 - 47424

  --1011100101000001    1011100101000010    1011100101000011    1011100101000100    1011100101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47425 - 47429

  --1011100101000110    1011100101000111    1011100101001000    1011100101001001    1011100101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47430 - 47434

  --1011100101001011    1011100101001100    1011100101001101    1011100101001110    1011100101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47435 - 47439

  --1011100101010000    1011100101010001    1011100101010010    1011100101010011    1011100101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47440 - 47444

  --1011100101010101    1011100101010110    1011100101010111    1011100101011000    1011100101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47445 - 47449

  --1011100101011010    1011100101011011    1011100101011100    1011100101011101    1011100101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47450 - 47454

  --1011100101011111    1011100101100000    1011100101100001    1011100101100010    1011100101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47455 - 47459

  --1011100101100100    1011100101100101    1011100101100110    1011100101100111    1011100101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47460 - 47464

  --1011100101101001    1011100101101010    1011100101101011    1011100101101100    1011100101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47465 - 47469

  --1011100101101110    1011100101101111    1011100101110000    1011100101110001    1011100101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47470 - 47474

  --1011100101110011    1011100101110100    1011100101110101    1011100101110110    1011100101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47475 - 47479

  --1011100101111000    1011100101111001    1011100101111010    1011100101111011    1011100101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47480 - 47484

  --1011100101111101    1011100101111110    1011100101111111    1011100110000000    1011100110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47485 - 47489

  --1011100110000010    1011100110000011    1011100110000100    1011100110000101    1011100110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47490 - 47494

  --1011100110000111    1011100110001000    1011100110001001    1011100110001010    1011100110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47495 - 47499

  --1011100110001100    1011100110001101    1011100110001110    1011100110001111    1011100110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47500 - 47504

  --1011100110010001    1011100110010010    1011100110010011    1011100110010100    1011100110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47505 - 47509

  --1011100110010110    1011100110010111    1011100110011000    1011100110011001    1011100110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47510 - 47514

  --1011100110011011    1011100110011100    1011100110011101    1011100110011110    1011100110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47515 - 47519

  --1011100110100000    1011100110100001    1011100110100010    1011100110100011    1011100110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47520 - 47524

  --1011100110100101    1011100110100110    1011100110100111    1011100110101000    1011100110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47525 - 47529

  --1011100110101010    1011100110101011    1011100110101100    1011100110101101    1011100110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47530 - 47534

  --1011100110101111    1011100110110000    1011100110110001    1011100110110010    1011100110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47535 - 47539

  --1011100110110100    1011100110110101    1011100110110110    1011100110110111    1011100110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47540 - 47544

  --1011100110111001    1011100110111010    1011100110111011    1011100110111100    1011100110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47545 - 47549

  --1011100110111110    1011100110111111    1011100111000000    1011100111000001    1011100111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47550 - 47554

  --1011100111000011    1011100111000100    1011100111000101    1011100111000110    1011100111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47555 - 47559

  --1011100111001000    1011100111001001    1011100111001010    1011100111001011    1011100111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47560 - 47564

  --1011100111001101    1011100111001110    1011100111001111    1011100111010000    1011100111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47565 - 47569

  --1011100111010010    1011100111010011    1011100111010100    1011100111010101    1011100111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47570 - 47574

  --1011100111010111    1011100111011000    1011100111011001    1011100111011010    1011100111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47575 - 47579

  --1011100111011100    1011100111011101    1011100111011110    1011100111011111    1011100111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47580 - 47584

  --1011100111100001    1011100111100010    1011100111100011    1011100111100100    1011100111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47585 - 47589

  --1011100111100110    1011100111100111    1011100111101000    1011100111101001    1011100111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47590 - 47594

  --1011100111101011    1011100111101100    1011100111101101    1011100111101110    1011100111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47595 - 47599

  --1011100111110000    1011100111110001    1011100111110010    1011100111110011    1011100111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47600 - 47604

  --1011100111110101    1011100111110110    1011100111110111    1011100111111000    1011100111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47605 - 47609

  --1011100111111010    1011100111111011    1011100111111100    1011100111111101    1011100111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47610 - 47614

  --1011100111111111    1011101000000000    1011101000000001    1011101000000010    1011101000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47615 - 47619

  --1011101000000100    1011101000000101    1011101000000110    1011101000000111    1011101000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47620 - 47624

  --1011101000001001    1011101000001010    1011101000001011    1011101000001100    1011101000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47625 - 47629

  --1011101000001110    1011101000001111    1011101000010000    1011101000010001    1011101000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47630 - 47634

  --1011101000010011    1011101000010100    1011101000010101    1011101000010110    1011101000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47635 - 47639

  --1011101000011000    1011101000011001    1011101000011010    1011101000011011    1011101000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47640 - 47644

  --1011101000011101    1011101000011110    1011101000011111    1011101000100000    1011101000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47645 - 47649

  --1011101000100010    1011101000100011    1011101000100100    1011101000100101    1011101000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47650 - 47654

  --1011101000100111    1011101000101000    1011101000101001    1011101000101010    1011101000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47655 - 47659

  --1011101000101100    1011101000101101    1011101000101110    1011101000101111    1011101000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47660 - 47664

  --1011101000110001    1011101000110010    1011101000110011    1011101000110100    1011101000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47665 - 47669

  --1011101000110110    1011101000110111    1011101000111000    1011101000111001    1011101000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47670 - 47674

  --1011101000111011    1011101000111100    1011101000111101    1011101000111110    1011101000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47675 - 47679

  --1011101001000000    1011101001000001    1011101001000010    1011101001000011    1011101001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47680 - 47684

  --1011101001000101    1011101001000110    1011101001000111    1011101001001000    1011101001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47685 - 47689

  --1011101001001010    1011101001001011    1011101001001100    1011101001001101    1011101001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47690 - 47694

  --1011101001001111    1011101001010000    1011101001010001    1011101001010010    1011101001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47695 - 47699

  --1011101001010100    1011101001010101    1011101001010110    1011101001010111    1011101001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47700 - 47704

  --1011101001011001    1011101001011010    1011101001011011    1011101001011100    1011101001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47705 - 47709

  --1011101001011110    1011101001011111    1011101001100000    1011101001100001    1011101001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47710 - 47714

  --1011101001100011    1011101001100100    1011101001100101    1011101001100110    1011101001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47715 - 47719

  --1011101001101000    1011101001101001    1011101001101010    1011101001101011    1011101001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47720 - 47724

  --1011101001101101    1011101001101110    1011101001101111    1011101001110000    1011101001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47725 - 47729

  --1011101001110010    1011101001110011    1011101001110100    1011101001110101    1011101001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47730 - 47734

  --1011101001110111    1011101001111000    1011101001111001    1011101001111010    1011101001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47735 - 47739

  --1011101001111100    1011101001111101    1011101001111110    1011101001111111    1011101010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47740 - 47744

  --1011101010000001    1011101010000010    1011101010000011    1011101010000100    1011101010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47745 - 47749

  --1011101010000110    1011101010000111    1011101010001000    1011101010001001    1011101010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47750 - 47754

  --1011101010001011    1011101010001100    1011101010001101    1011101010001110    1011101010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47755 - 47759

  --1011101010010000    1011101010010001    1011101010010010    1011101010010011    1011101010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47760 - 47764

  --1011101010010101    1011101010010110    1011101010010111    1011101010011000    1011101010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47765 - 47769

  --1011101010011010    1011101010011011    1011101010011100    1011101010011101    1011101010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47770 - 47774

  --1011101010011111    1011101010100000    1011101010100001    1011101010100010    1011101010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47775 - 47779

  --1011101010100100    1011101010100101    1011101010100110    1011101010100111    1011101010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47780 - 47784

  --1011101010101001    1011101010101010    1011101010101011    1011101010101100    1011101010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47785 - 47789

  --1011101010101110    1011101010101111    1011101010110000    1011101010110001    1011101010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47790 - 47794

  --1011101010110011    1011101010110100    1011101010110101    1011101010110110    1011101010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47795 - 47799

  --1011101010111000    1011101010111001    1011101010111010    1011101010111011    1011101010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47800 - 47804

  --1011101010111101    1011101010111110    1011101010111111    1011101011000000    1011101011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47805 - 47809

  --1011101011000010    1011101011000011    1011101011000100    1011101011000101    1011101011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47810 - 47814

  --1011101011000111    1011101011001000    1011101011001001    1011101011001010    1011101011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47815 - 47819

  --1011101011001100    1011101011001101    1011101011001110    1011101011001111    1011101011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47820 - 47824

  --1011101011010001    1011101011010010    1011101011010011    1011101011010100    1011101011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47825 - 47829

  --1011101011010110    1011101011010111    1011101011011000    1011101011011001    1011101011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47830 - 47834

  --1011101011011011    1011101011011100    1011101011011101    1011101011011110    1011101011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47835 - 47839

  --1011101011100000    1011101011100001    1011101011100010    1011101011100011    1011101011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47840 - 47844

  --1011101011100101    1011101011100110    1011101011100111    1011101011101000    1011101011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47845 - 47849

  --1011101011101010    1011101011101011    1011101011101100    1011101011101101    1011101011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47850 - 47854

  --1011101011101111    1011101011110000    1011101011110001    1011101011110010    1011101011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47855 - 47859

  --1011101011110100    1011101011110101    1011101011110110    1011101011110111    1011101011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47860 - 47864

  --1011101011111001    1011101011111010    1011101011111011    1011101011111100    1011101011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47865 - 47869

  --1011101011111110    1011101011111111    1011101100000000    1011101100000001    1011101100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47870 - 47874

  --1011101100000011    1011101100000100    1011101100000101    1011101100000110    1011101100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47875 - 47879

  --1011101100001000    1011101100001001    1011101100001010    1011101100001011    1011101100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47880 - 47884

  --1011101100001101    1011101100001110    1011101100001111    1011101100010000    1011101100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47885 - 47889

  --1011101100010010    1011101100010011    1011101100010100    1011101100010101    1011101100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47890 - 47894

  --1011101100010111    1011101100011000    1011101100011001    1011101100011010    1011101100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47895 - 47899

  --1011101100011100    1011101100011101    1011101100011110    1011101100011111    1011101100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47900 - 47904

  --1011101100100001    1011101100100010    1011101100100011    1011101100100100    1011101100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47905 - 47909

  --1011101100100110    1011101100100111    1011101100101000    1011101100101001    1011101100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47910 - 47914

  --1011101100101011    1011101100101100    1011101100101101    1011101100101110    1011101100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47915 - 47919

  --1011101100110000    1011101100110001    1011101100110010    1011101100110011    1011101100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47920 - 47924

  --1011101100110101    1011101100110110    1011101100110111    1011101100111000    1011101100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47925 - 47929

  --1011101100111010    1011101100111011    1011101100111100    1011101100111101    1011101100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47930 - 47934

  --1011101100111111    1011101101000000    1011101101000001    1011101101000010    1011101101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47935 - 47939

  --1011101101000100    1011101101000101    1011101101000110    1011101101000111    1011101101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47940 - 47944

  --1011101101001001    1011101101001010    1011101101001011    1011101101001100    1011101101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47945 - 47949

  --1011101101001110    1011101101001111    1011101101010000    1011101101010001    1011101101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47950 - 47954

  --1011101101010011    1011101101010100    1011101101010101    1011101101010110    1011101101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47955 - 47959

  --1011101101011000    1011101101011001    1011101101011010    1011101101011011    1011101101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47960 - 47964

  --1011101101011101    1011101101011110    1011101101011111    1011101101100000    1011101101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47965 - 47969

  --1011101101100010    1011101101100011    1011101101100100    1011101101100101    1011101101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47970 - 47974

  --1011101101100111    1011101101101000    1011101101101001    1011101101101010    1011101101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47975 - 47979

  --1011101101101100    1011101101101101    1011101101101110    1011101101101111    1011101101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47980 - 47984

  --1011101101110001    1011101101110010    1011101101110011    1011101101110100    1011101101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47985 - 47989

  --1011101101110110    1011101101110111    1011101101111000    1011101101111001    1011101101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47990 - 47994

  --1011101101111011    1011101101111100    1011101101111101    1011101101111110    1011101101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 47995 - 47999

  --1011101110000000    1011101110000001    1011101110000010    1011101110000011    1011101110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48000 - 48004

  --1011101110000101    1011101110000110    1011101110000111    1011101110001000    1011101110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48005 - 48009

  --1011101110001010    1011101110001011    1011101110001100    1011101110001101    1011101110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48010 - 48014

  --1011101110001111    1011101110010000    1011101110010001    1011101110010010    1011101110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48015 - 48019

  --1011101110010100    1011101110010101    1011101110010110    1011101110010111    1011101110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48020 - 48024

  --1011101110011001    1011101110011010    1011101110011011    1011101110011100    1011101110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48025 - 48029

  --1011101110011110    1011101110011111    1011101110100000    1011101110100001    1011101110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48030 - 48034

  --1011101110100011    1011101110100100    1011101110100101    1011101110100110    1011101110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48035 - 48039

  --1011101110101000    1011101110101001    1011101110101010    1011101110101011    1011101110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48040 - 48044

  --1011101110101101    1011101110101110    1011101110101111    1011101110110000    1011101110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48045 - 48049

  --1011101110110010    1011101110110011    1011101110110100    1011101110110101    1011101110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48050 - 48054

  --1011101110110111    1011101110111000    1011101110111001    1011101110111010    1011101110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48055 - 48059

  --1011101110111100    1011101110111101    1011101110111110    1011101110111111    1011101111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48060 - 48064

  --1011101111000001    1011101111000010    1011101111000011    1011101111000100    1011101111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48065 - 48069

  --1011101111000110    1011101111000111    1011101111001000    1011101111001001    1011101111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48070 - 48074

  --1011101111001011    1011101111001100    1011101111001101    1011101111001110    1011101111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48075 - 48079

  --1011101111010000    1011101111010001    1011101111010010    1011101111010011    1011101111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48080 - 48084

  --1011101111010101    1011101111010110    1011101111010111    1011101111011000    1011101111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48085 - 48089

  --1011101111011010    1011101111011011    1011101111011100    1011101111011101    1011101111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48090 - 48094

  --1011101111011111    1011101111100000    1011101111100001    1011101111100010    1011101111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48095 - 48099

  --1011101111100100    1011101111100101    1011101111100110    1011101111100111    1011101111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48100 - 48104

  --1011101111101001    1011101111101010    1011101111101011    1011101111101100    1011101111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48105 - 48109

  --1011101111101110    1011101111101111    1011101111110000    1011101111110001    1011101111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48110 - 48114

  --1011101111110011    1011101111110100    1011101111110101    1011101111110110    1011101111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48115 - 48119

  --1011101111111000    1011101111111001    1011101111111010    1011101111111011    1011101111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48120 - 48124

  --1011101111111101    1011101111111110    1011101111111111    1011110000000000    1011110000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48125 - 48129

  --1011110000000010    1011110000000011    1011110000000100    1011110000000101    1011110000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48130 - 48134

  --1011110000000111    1011110000001000    1011110000001001    1011110000001010    1011110000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48135 - 48139

  --1011110000001100    1011110000001101    1011110000001110    1011110000001111    1011110000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48140 - 48144

  --1011110000010001    1011110000010010    1011110000010011    1011110000010100    1011110000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48145 - 48149

  --1011110000010110    1011110000010111    1011110000011000    1011110000011001    1011110000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48150 - 48154

  --1011110000011011    1011110000011100    1011110000011101    1011110000011110    1011110000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48155 - 48159

  --1011110000100000    1011110000100001    1011110000100010    1011110000100011    1011110000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48160 - 48164

  --1011110000100101    1011110000100110    1011110000100111    1011110000101000    1011110000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48165 - 48169

  --1011110000101010    1011110000101011    1011110000101100    1011110000101101    1011110000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48170 - 48174

  --1011110000101111    1011110000110000    1011110000110001    1011110000110010    1011110000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48175 - 48179

  --1011110000110100    1011110000110101    1011110000110110    1011110000110111    1011110000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48180 - 48184

  --1011110000111001    1011110000111010    1011110000111011    1011110000111100    1011110000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48185 - 48189

  --1011110000111110    1011110000111111    1011110001000000    1011110001000001    1011110001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48190 - 48194

  --1011110001000011    1011110001000100    1011110001000101    1011110001000110    1011110001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48195 - 48199

  --1011110001001000    1011110001001001    1011110001001010    1011110001001011    1011110001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48200 - 48204

  --1011110001001101    1011110001001110    1011110001001111    1011110001010000    1011110001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48205 - 48209

  --1011110001010010    1011110001010011    1011110001010100    1011110001010101    1011110001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48210 - 48214

  --1011110001010111    1011110001011000    1011110001011001    1011110001011010    1011110001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48215 - 48219

  --1011110001011100    1011110001011101    1011110001011110    1011110001011111    1011110001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48220 - 48224

  --1011110001100001    1011110001100010    1011110001100011    1011110001100100    1011110001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48225 - 48229

  --1011110001100110    1011110001100111    1011110001101000    1011110001101001    1011110001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48230 - 48234

  --1011110001101011    1011110001101100    1011110001101101    1011110001101110    1011110001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48235 - 48239

  --1011110001110000    1011110001110001    1011110001110010    1011110001110011    1011110001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48240 - 48244

  --1011110001110101    1011110001110110    1011110001110111    1011110001111000    1011110001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48245 - 48249

  --1011110001111010    1011110001111011    1011110001111100    1011110001111101    1011110001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48250 - 48254

  --1011110001111111    1011110010000000    1011110010000001    1011110010000010    1011110010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48255 - 48259

  --1011110010000100    1011110010000101    1011110010000110    1011110010000111    1011110010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48260 - 48264

  --1011110010001001    1011110010001010    1011110010001011    1011110010001100    1011110010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48265 - 48269

  --1011110010001110    1011110010001111    1011110010010000    1011110010010001    1011110010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48270 - 48274

  --1011110010010011    1011110010010100    1011110010010101    1011110010010110    1011110010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48275 - 48279

  --1011110010011000    1011110010011001    1011110010011010    1011110010011011    1011110010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48280 - 48284

  --1011110010011101    1011110010011110    1011110010011111    1011110010100000    1011110010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48285 - 48289

  --1011110010100010    1011110010100011    1011110010100100    1011110010100101    1011110010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48290 - 48294

  --1011110010100111    1011110010101000    1011110010101001    1011110010101010    1011110010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48295 - 48299

  --1011110010101100    1011110010101101    1011110010101110    1011110010101111    1011110010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48300 - 48304

  --1011110010110001    1011110010110010    1011110010110011    1011110010110100    1011110010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48305 - 48309

  --1011110010110110    1011110010110111    1011110010111000    1011110010111001    1011110010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48310 - 48314

  --1011110010111011    1011110010111100    1011110010111101    1011110010111110    1011110010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48315 - 48319

  --1011110011000000    1011110011000001    1011110011000010    1011110011000011    1011110011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48320 - 48324

  --1011110011000101    1011110011000110    1011110011000111    1011110011001000    1011110011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48325 - 48329

  --1011110011001010    1011110011001011    1011110011001100    1011110011001101    1011110011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48330 - 48334

  --1011110011001111    1011110011010000    1011110011010001    1011110011010010    1011110011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48335 - 48339

  --1011110011010100    1011110011010101    1011110011010110    1011110011010111    1011110011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48340 - 48344

  --1011110011011001    1011110011011010    1011110011011011    1011110011011100    1011110011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48345 - 48349

  --1011110011011110    1011110011011111    1011110011100000    1011110011100001    1011110011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48350 - 48354

  --1011110011100011    1011110011100100    1011110011100101    1011110011100110    1011110011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48355 - 48359

  --1011110011101000    1011110011101001    1011110011101010    1011110011101011    1011110011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48360 - 48364

  --1011110011101101    1011110011101110    1011110011101111    1011110011110000    1011110011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48365 - 48369

  --1011110011110010    1011110011110011    1011110011110100    1011110011110101    1011110011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48370 - 48374

  --1011110011110111    1011110011111000    1011110011111001    1011110011111010    1011110011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48375 - 48379

  --1011110011111100    1011110011111101    1011110011111110    1011110011111111    1011110100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48380 - 48384

  --1011110100000001    1011110100000010    1011110100000011    1011110100000100    1011110100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48385 - 48389

  --1011110100000110    1011110100000111    1011110100001000    1011110100001001    1011110100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48390 - 48394

  --1011110100001011    1011110100001100    1011110100001101    1011110100001110    1011110100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48395 - 48399

  --1011110100010000    1011110100010001    1011110100010010    1011110100010011    1011110100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48400 - 48404

  --1011110100010101    1011110100010110    1011110100010111    1011110100011000    1011110100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48405 - 48409

  --1011110100011010    1011110100011011    1011110100011100    1011110100011101    1011110100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48410 - 48414

  --1011110100011111    1011110100100000    1011110100100001    1011110100100010    1011110100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48415 - 48419

  --1011110100100100    1011110100100101    1011110100100110    1011110100100111    1011110100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48420 - 48424

  --1011110100101001    1011110100101010    1011110100101011    1011110100101100    1011110100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48425 - 48429

  --1011110100101110    1011110100101111    1011110100110000    1011110100110001    1011110100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48430 - 48434

  --1011110100110011    1011110100110100    1011110100110101    1011110100110110    1011110100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48435 - 48439

  --1011110100111000    1011110100111001    1011110100111010    1011110100111011    1011110100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48440 - 48444

  --1011110100111101    1011110100111110    1011110100111111    1011110101000000    1011110101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48445 - 48449

  --1011110101000010    1011110101000011    1011110101000100    1011110101000101    1011110101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48450 - 48454

  --1011110101000111    1011110101001000    1011110101001001    1011110101001010    1011110101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48455 - 48459

  --1011110101001100    1011110101001101    1011110101001110    1011110101001111    1011110101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48460 - 48464

  --1011110101010001    1011110101010010    1011110101010011    1011110101010100    1011110101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48465 - 48469

  --1011110101010110    1011110101010111    1011110101011000    1011110101011001    1011110101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48470 - 48474

  --1011110101011011    1011110101011100    1011110101011101    1011110101011110    1011110101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48475 - 48479

  --1011110101100000    1011110101100001    1011110101100010    1011110101100011    1011110101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48480 - 48484

  --1011110101100101    1011110101100110    1011110101100111    1011110101101000    1011110101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48485 - 48489

  --1011110101101010    1011110101101011    1011110101101100    1011110101101101    1011110101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48490 - 48494

  --1011110101101111    1011110101110000    1011110101110001    1011110101110010    1011110101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48495 - 48499

  --1011110101110100    1011110101110101    1011110101110110    1011110101110111    1011110101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48500 - 48504

  --1011110101111001    1011110101111010    1011110101111011    1011110101111100    1011110101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48505 - 48509

  --1011110101111110    1011110101111111    1011110110000000    1011110110000001    1011110110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48510 - 48514

  --1011110110000011    1011110110000100    1011110110000101    1011110110000110    1011110110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48515 - 48519

  --1011110110001000    1011110110001001    1011110110001010    1011110110001011    1011110110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48520 - 48524

  --1011110110001101    1011110110001110    1011110110001111    1011110110010000    1011110110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48525 - 48529

  --1011110110010010    1011110110010011    1011110110010100    1011110110010101    1011110110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48530 - 48534

  --1011110110010111    1011110110011000    1011110110011001    1011110110011010    1011110110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48535 - 48539

  --1011110110011100    1011110110011101    1011110110011110    1011110110011111    1011110110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48540 - 48544

  --1011110110100001    1011110110100010    1011110110100011    1011110110100100    1011110110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48545 - 48549

  --1011110110100110    1011110110100111    1011110110101000    1011110110101001    1011110110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48550 - 48554

  --1011110110101011    1011110110101100    1011110110101101    1011110110101110    1011110110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48555 - 48559

  --1011110110110000    1011110110110001    1011110110110010    1011110110110011    1011110110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48560 - 48564

  --1011110110110101    1011110110110110    1011110110110111    1011110110111000    1011110110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48565 - 48569

  --1011110110111010    1011110110111011    1011110110111100    1011110110111101    1011110110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48570 - 48574

  --1011110110111111    1011110111000000    1011110111000001    1011110111000010    1011110111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48575 - 48579

  --1011110111000100    1011110111000101    1011110111000110    1011110111000111    1011110111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48580 - 48584

  --1011110111001001    1011110111001010    1011110111001011    1011110111001100    1011110111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48585 - 48589

  --1011110111001110    1011110111001111    1011110111010000    1011110111010001    1011110111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48590 - 48594

  --1011110111010011    1011110111010100    1011110111010101    1011110111010110    1011110111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48595 - 48599

  --1011110111011000    1011110111011001    1011110111011010    1011110111011011    1011110111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48600 - 48604

  --1011110111011101    1011110111011110    1011110111011111    1011110111100000    1011110111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48605 - 48609

  --1011110111100010    1011110111100011    1011110111100100    1011110111100101    1011110111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48610 - 48614

  --1011110111100111    1011110111101000    1011110111101001    1011110111101010    1011110111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48615 - 48619

  --1011110111101100    1011110111101101    1011110111101110    1011110111101111    1011110111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48620 - 48624

  --1011110111110001    1011110111110010    1011110111110011    1011110111110100    1011110111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48625 - 48629

  --1011110111110110    1011110111110111    1011110111111000    1011110111111001    1011110111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48630 - 48634

  --1011110111111011    1011110111111100    1011110111111101    1011110111111110    1011110111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48635 - 48639

  --1011111000000000    1011111000000001    1011111000000010    1011111000000011    1011111000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48640 - 48644

  --1011111000000101    1011111000000110    1011111000000111    1011111000001000    1011111000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48645 - 48649

  --1011111000001010    1011111000001011    1011111000001100    1011111000001101    1011111000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48650 - 48654

  --1011111000001111    1011111000010000    1011111000010001    1011111000010010    1011111000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48655 - 48659

  --1011111000010100    1011111000010101    1011111000010110    1011111000010111    1011111000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48660 - 48664

  --1011111000011001    1011111000011010    1011111000011011    1011111000011100    1011111000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48665 - 48669

  --1011111000011110    1011111000011111    1011111000100000    1011111000100001    1011111000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48670 - 48674

  --1011111000100011    1011111000100100    1011111000100101    1011111000100110    1011111000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48675 - 48679

  --1011111000101000    1011111000101001    1011111000101010    1011111000101011    1011111000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48680 - 48684

  --1011111000101101    1011111000101110    1011111000101111    1011111000110000    1011111000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48685 - 48689

  --1011111000110010    1011111000110011    1011111000110100    1011111000110101    1011111000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48690 - 48694

  --1011111000110111    1011111000111000    1011111000111001    1011111000111010    1011111000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48695 - 48699

  --1011111000111100    1011111000111101    1011111000111110    1011111000111111    1011111001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48700 - 48704

  --1011111001000001    1011111001000010    1011111001000011    1011111001000100    1011111001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48705 - 48709

  --1011111001000110    1011111001000111    1011111001001000    1011111001001001    1011111001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48710 - 48714

  --1011111001001011    1011111001001100    1011111001001101    1011111001001110    1011111001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48715 - 48719

  --1011111001010000    1011111001010001    1011111001010010    1011111001010011    1011111001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48720 - 48724

  --1011111001010101    1011111001010110    1011111001010111    1011111001011000    1011111001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48725 - 48729

  --1011111001011010    1011111001011011    1011111001011100    1011111001011101    1011111001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48730 - 48734

  --1011111001011111    1011111001100000    1011111001100001    1011111001100010    1011111001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48735 - 48739

  --1011111001100100    1011111001100101    1011111001100110    1011111001100111    1011111001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48740 - 48744

  --1011111001101001    1011111001101010    1011111001101011    1011111001101100    1011111001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48745 - 48749

  --1011111001101110    1011111001101111    1011111001110000    1011111001110001    1011111001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48750 - 48754

  --1011111001110011    1011111001110100    1011111001110101    1011111001110110    1011111001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48755 - 48759

  --1011111001111000    1011111001111001    1011111001111010    1011111001111011    1011111001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48760 - 48764

  --1011111001111101    1011111001111110    1011111001111111    1011111010000000    1011111010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48765 - 48769

  --1011111010000010    1011111010000011    1011111010000100    1011111010000101    1011111010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48770 - 48774

  --1011111010000111    1011111010001000    1011111010001001    1011111010001010    1011111010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48775 - 48779

  --1011111010001100    1011111010001101    1011111010001110    1011111010001111    1011111010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48780 - 48784

  --1011111010010001    1011111010010010    1011111010010011    1011111010010100    1011111010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48785 - 48789

  --1011111010010110    1011111010010111    1011111010011000    1011111010011001    1011111010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48790 - 48794

  --1011111010011011    1011111010011100    1011111010011101    1011111010011110    1011111010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48795 - 48799

  --1011111010100000    1011111010100001    1011111010100010    1011111010100011    1011111010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48800 - 48804

  --1011111010100101    1011111010100110    1011111010100111    1011111010101000    1011111010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48805 - 48809

  --1011111010101010    1011111010101011    1011111010101100    1011111010101101    1011111010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48810 - 48814

  --1011111010101111    1011111010110000    1011111010110001    1011111010110010    1011111010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48815 - 48819

  --1011111010110100    1011111010110101    1011111010110110    1011111010110111    1011111010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48820 - 48824

  --1011111010111001    1011111010111010    1011111010111011    1011111010111100    1011111010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48825 - 48829

  --1011111010111110    1011111010111111    1011111011000000    1011111011000001    1011111011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48830 - 48834

  --1011111011000011    1011111011000100    1011111011000101    1011111011000110    1011111011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48835 - 48839

  --1011111011001000    1011111011001001    1011111011001010    1011111011001011    1011111011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48840 - 48844

  --1011111011001101    1011111011001110    1011111011001111    1011111011010000    1011111011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48845 - 48849

  --1011111011010010    1011111011010011    1011111011010100    1011111011010101    1011111011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48850 - 48854

  --1011111011010111    1011111011011000    1011111011011001    1011111011011010    1011111011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48855 - 48859

  --1011111011011100    1011111011011101    1011111011011110    1011111011011111    1011111011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48860 - 48864

  --1011111011100001    1011111011100010    1011111011100011    1011111011100100    1011111011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48865 - 48869

  --1011111011100110    1011111011100111    1011111011101000    1011111011101001    1011111011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48870 - 48874

  --1011111011101011    1011111011101100    1011111011101101    1011111011101110    1011111011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48875 - 48879

  --1011111011110000    1011111011110001    1011111011110010    1011111011110011    1011111011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48880 - 48884

  --1011111011110101    1011111011110110    1011111011110111    1011111011111000    1011111011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48885 - 48889

  --1011111011111010    1011111011111011    1011111011111100    1011111011111101    1011111011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48890 - 48894

  --1011111011111111    1011111100000000    1011111100000001    1011111100000010    1011111100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48895 - 48899

  --1011111100000100    1011111100000101    1011111100000110    1011111100000111    1011111100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48900 - 48904

  --1011111100001001    1011111100001010    1011111100001011    1011111100001100    1011111100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48905 - 48909

  --1011111100001110    1011111100001111    1011111100010000    1011111100010001    1011111100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48910 - 48914

  --1011111100010011    1011111100010100    1011111100010101    1011111100010110    1011111100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48915 - 48919

  --1011111100011000    1011111100011001    1011111100011010    1011111100011011    1011111100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48920 - 48924

  --1011111100011101    1011111100011110    1011111100011111    1011111100100000    1011111100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48925 - 48929

  --1011111100100010    1011111100100011    1011111100100100    1011111100100101    1011111100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48930 - 48934

  --1011111100100111    1011111100101000    1011111100101001    1011111100101010    1011111100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48935 - 48939

  --1011111100101100    1011111100101101    1011111100101110    1011111100101111    1011111100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48940 - 48944

  --1011111100110001    1011111100110010    1011111100110011    1011111100110100    1011111100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48945 - 48949

  --1011111100110110    1011111100110111    1011111100111000    1011111100111001    1011111100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48950 - 48954

  --1011111100111011    1011111100111100    1011111100111101    1011111100111110    1011111100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48955 - 48959

  --1011111101000000    1011111101000001    1011111101000010    1011111101000011    1011111101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48960 - 48964

  --1011111101000101    1011111101000110    1011111101000111    1011111101001000    1011111101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48965 - 48969

  --1011111101001010    1011111101001011    1011111101001100    1011111101001101    1011111101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48970 - 48974

  --1011111101001111    1011111101010000    1011111101010001    1011111101010010    1011111101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48975 - 48979

  --1011111101010100    1011111101010101    1011111101010110    1011111101010111    1011111101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48980 - 48984

  --1011111101011001    1011111101011010    1011111101011011    1011111101011100    1011111101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48985 - 48989

  --1011111101011110    1011111101011111    1011111101100000    1011111101100001    1011111101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48990 - 48994

  --1011111101100011    1011111101100100    1011111101100101    1011111101100110    1011111101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 48995 - 48999

  --1011111101101000    1011111101101001    1011111101101010    1011111101101011    1011111101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49000 - 49004

  --1011111101101101    1011111101101110    1011111101101111    1011111101110000    1011111101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49005 - 49009

  --1011111101110010    1011111101110011    1011111101110100    1011111101110101    1011111101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49010 - 49014

  --1011111101110111    1011111101111000    1011111101111001    1011111101111010    1011111101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49015 - 49019

  --1011111101111100    1011111101111101    1011111101111110    1011111101111111    1011111110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49020 - 49024

  --1011111110000001    1011111110000010    1011111110000011    1011111110000100    1011111110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49025 - 49029

  --1011111110000110    1011111110000111    1011111110001000    1011111110001001    1011111110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49030 - 49034

  --1011111110001011    1011111110001100    1011111110001101    1011111110001110    1011111110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49035 - 49039

  --1011111110010000    1011111110010001    1011111110010010    1011111110010011    1011111110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49040 - 49044

  --1011111110010101    1011111110010110    1011111110010111    1011111110011000    1011111110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49045 - 49049

  --1011111110011010    1011111110011011    1011111110011100    1011111110011101    1011111110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49050 - 49054

  --1011111110011111    1011111110100000    1011111110100001    1011111110100010    1011111110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49055 - 49059

  --1011111110100100    1011111110100101    1011111110100110    1011111110100111    1011111110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49060 - 49064

  --1011111110101001    1011111110101010    1011111110101011    1011111110101100    1011111110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49065 - 49069

  --1011111110101110    1011111110101111    1011111110110000    1011111110110001    1011111110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49070 - 49074

  --1011111110110011    1011111110110100    1011111110110101    1011111110110110    1011111110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49075 - 49079

  --1011111110111000    1011111110111001    1011111110111010    1011111110111011    1011111110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49080 - 49084

  --1011111110111101    1011111110111110    1011111110111111    1011111111000000    1011111111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49085 - 49089

  --1011111111000010    1011111111000011    1011111111000100    1011111111000101    1011111111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49090 - 49094

  --1011111111000111    1011111111001000    1011111111001001    1011111111001010    1011111111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49095 - 49099

  --1011111111001100    1011111111001101    1011111111001110    1011111111001111    1011111111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49100 - 49104

  --1011111111010001    1011111111010010    1011111111010011    1011111111010100    1011111111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49105 - 49109

  --1011111111010110    1011111111010111    1011111111011000    1011111111011001    1011111111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49110 - 49114

  --1011111111011011    1011111111011100    1011111111011101    1011111111011110    1011111111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49115 - 49119

  --1011111111100000    1011111111100001    1011111111100010    1011111111100011    1011111111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49120 - 49124

  --1011111111100101    1011111111100110    1011111111100111    1011111111101000    1011111111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49125 - 49129

  --1011111111101010    1011111111101011    1011111111101100    1011111111101101    1011111111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49130 - 49134

  --1011111111101111    1011111111110000    1011111111110001    1011111111110010    1011111111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49135 - 49139

  --1011111111110100    1011111111110101    1011111111110110    1011111111110111    1011111111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49140 - 49144

  --1011111111111001    1011111111111010    1011111111111011    1011111111111100    1011111111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49145 - 49149

  --1011111111111110    1011111111111111    1100000000000000    1100000000000001    1100000000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49150 - 49154

  --1100000000000011    1100000000000100    1100000000000101    1100000000000110    1100000000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49155 - 49159

  --1100000000001000    1100000000001001    1100000000001010    1100000000001011    1100000000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49160 - 49164

  --1100000000001101    1100000000001110    1100000000001111    1100000000010000    1100000000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49165 - 49169

  --1100000000010010    1100000000010011    1100000000010100    1100000000010101    1100000000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49170 - 49174

  --1100000000010111    1100000000011000    1100000000011001    1100000000011010    1100000000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49175 - 49179

  --1100000000011100    1100000000011101    1100000000011110    1100000000011111    1100000000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49180 - 49184

  --1100000000100001    1100000000100010    1100000000100011    1100000000100100    1100000000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49185 - 49189

  --1100000000100110    1100000000100111    1100000000101000    1100000000101001    1100000000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49190 - 49194

  --1100000000101011    1100000000101100    1100000000101101    1100000000101110    1100000000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49195 - 49199

  --1100000000110000    1100000000110001    1100000000110010    1100000000110011    1100000000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49200 - 49204

  --1100000000110101    1100000000110110    1100000000110111    1100000000111000    1100000000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49205 - 49209

  --1100000000111010    1100000000111011    1100000000111100    1100000000111101    1100000000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49210 - 49214

  --1100000000111111    1100000001000000    1100000001000001    1100000001000010    1100000001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49215 - 49219

  --1100000001000100    1100000001000101    1100000001000110    1100000001000111    1100000001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49220 - 49224

  --1100000001001001    1100000001001010    1100000001001011    1100000001001100    1100000001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49225 - 49229

  --1100000001001110    1100000001001111    1100000001010000    1100000001010001    1100000001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49230 - 49234

  --1100000001010011    1100000001010100    1100000001010101    1100000001010110    1100000001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49235 - 49239

  --1100000001011000    1100000001011001    1100000001011010    1100000001011011    1100000001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49240 - 49244

  --1100000001011101    1100000001011110    1100000001011111    1100000001100000    1100000001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49245 - 49249

  --1100000001100010    1100000001100011    1100000001100100    1100000001100101    1100000001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49250 - 49254

  --1100000001100111    1100000001101000    1100000001101001    1100000001101010    1100000001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49255 - 49259

  --1100000001101100    1100000001101101    1100000001101110    1100000001101111    1100000001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49260 - 49264

  --1100000001110001    1100000001110010    1100000001110011    1100000001110100    1100000001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49265 - 49269

  --1100000001110110    1100000001110111    1100000001111000    1100000001111001    1100000001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49270 - 49274

  --1100000001111011    1100000001111100    1100000001111101    1100000001111110    1100000001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49275 - 49279

  --1100000010000000    1100000010000001    1100000010000010    1100000010000011    1100000010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49280 - 49284

  --1100000010000101    1100000010000110    1100000010000111    1100000010001000    1100000010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49285 - 49289

  --1100000010001010    1100000010001011    1100000010001100    1100000010001101    1100000010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49290 - 49294

  --1100000010001111    1100000010010000    1100000010010001    1100000010010010    1100000010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49295 - 49299

  --1100000010010100    1100000010010101    1100000010010110    1100000010010111    1100000010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49300 - 49304

  --1100000010011001    1100000010011010    1100000010011011    1100000010011100    1100000010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49305 - 49309

  --1100000010011110    1100000010011111    1100000010100000    1100000010100001    1100000010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49310 - 49314

  --1100000010100011    1100000010100100    1100000010100101    1100000010100110    1100000010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49315 - 49319

  --1100000010101000    1100000010101001    1100000010101010    1100000010101011    1100000010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49320 - 49324

  --1100000010101101    1100000010101110    1100000010101111    1100000010110000    1100000010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49325 - 49329

  --1100000010110010    1100000010110011    1100000010110100    1100000010110101    1100000010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49330 - 49334

  --1100000010110111    1100000010111000    1100000010111001    1100000010111010    1100000010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49335 - 49339

  --1100000010111100    1100000010111101    1100000010111110    1100000010111111    1100000011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49340 - 49344

  --1100000011000001    1100000011000010    1100000011000011    1100000011000100    1100000011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49345 - 49349

  --1100000011000110    1100000011000111    1100000011001000    1100000011001001    1100000011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49350 - 49354

  --1100000011001011    1100000011001100    1100000011001101    1100000011001110    1100000011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49355 - 49359

  --1100000011010000    1100000011010001    1100000011010010    1100000011010011    1100000011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49360 - 49364

  --1100000011010101    1100000011010110    1100000011010111    1100000011011000    1100000011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49365 - 49369

  --1100000011011010    1100000011011011    1100000011011100    1100000011011101    1100000011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49370 - 49374

  --1100000011011111    1100000011100000    1100000011100001    1100000011100010    1100000011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49375 - 49379

  --1100000011100100    1100000011100101    1100000011100110    1100000011100111    1100000011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49380 - 49384

  --1100000011101001    1100000011101010    1100000011101011    1100000011101100    1100000011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49385 - 49389

  --1100000011101110    1100000011101111    1100000011110000    1100000011110001    1100000011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49390 - 49394

  --1100000011110011    1100000011110100    1100000011110101    1100000011110110    1100000011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49395 - 49399

  --1100000011111000    1100000011111001    1100000011111010    1100000011111011    1100000011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49400 - 49404

  --1100000011111101    1100000011111110    1100000011111111    1100000100000000    1100000100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49405 - 49409

  --1100000100000010    1100000100000011    1100000100000100    1100000100000101    1100000100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49410 - 49414

  --1100000100000111    1100000100001000    1100000100001001    1100000100001010    1100000100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49415 - 49419

  --1100000100001100    1100000100001101    1100000100001110    1100000100001111    1100000100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49420 - 49424

  --1100000100010001    1100000100010010    1100000100010011    1100000100010100    1100000100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49425 - 49429

  --1100000100010110    1100000100010111    1100000100011000    1100000100011001    1100000100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49430 - 49434

  --1100000100011011    1100000100011100    1100000100011101    1100000100011110    1100000100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49435 - 49439

  --1100000100100000    1100000100100001    1100000100100010    1100000100100011    1100000100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49440 - 49444

  --1100000100100101    1100000100100110    1100000100100111    1100000100101000    1100000100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49445 - 49449

  --1100000100101010    1100000100101011    1100000100101100    1100000100101101    1100000100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49450 - 49454

  --1100000100101111    1100000100110000    1100000100110001    1100000100110010    1100000100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49455 - 49459

  --1100000100110100    1100000100110101    1100000100110110    1100000100110111    1100000100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49460 - 49464

  --1100000100111001    1100000100111010    1100000100111011    1100000100111100    1100000100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49465 - 49469

  --1100000100111110    1100000100111111    1100000101000000    1100000101000001    1100000101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49470 - 49474

  --1100000101000011    1100000101000100    1100000101000101    1100000101000110    1100000101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49475 - 49479

  --1100000101001000    1100000101001001    1100000101001010    1100000101001011    1100000101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49480 - 49484

  --1100000101001101    1100000101001110    1100000101001111    1100000101010000    1100000101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49485 - 49489

  --1100000101010010    1100000101010011    1100000101010100    1100000101010101    1100000101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49490 - 49494

  --1100000101010111    1100000101011000    1100000101011001    1100000101011010    1100000101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49495 - 49499

  --1100000101011100    1100000101011101    1100000101011110    1100000101011111    1100000101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49500 - 49504

  --1100000101100001    1100000101100010    1100000101100011    1100000101100100    1100000101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49505 - 49509

  --1100000101100110    1100000101100111    1100000101101000    1100000101101001    1100000101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49510 - 49514

  --1100000101101011    1100000101101100    1100000101101101    1100000101101110    1100000101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49515 - 49519

  --1100000101110000    1100000101110001    1100000101110010    1100000101110011    1100000101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49520 - 49524

  --1100000101110101    1100000101110110    1100000101110111    1100000101111000    1100000101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49525 - 49529

  --1100000101111010    1100000101111011    1100000101111100    1100000101111101    1100000101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49530 - 49534

  --1100000101111111    1100000110000000    1100000110000001    1100000110000010    1100000110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49535 - 49539

  --1100000110000100    1100000110000101    1100000110000110    1100000110000111    1100000110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49540 - 49544

  --1100000110001001    1100000110001010    1100000110001011    1100000110001100    1100000110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49545 - 49549

  --1100000110001110    1100000110001111    1100000110010000    1100000110010001    1100000110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49550 - 49554

  --1100000110010011    1100000110010100    1100000110010101    1100000110010110    1100000110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49555 - 49559

  --1100000110011000    1100000110011001    1100000110011010    1100000110011011    1100000110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49560 - 49564

  --1100000110011101    1100000110011110    1100000110011111    1100000110100000    1100000110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49565 - 49569

  --1100000110100010    1100000110100011    1100000110100100    1100000110100101    1100000110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49570 - 49574

  --1100000110100111    1100000110101000    1100000110101001    1100000110101010    1100000110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49575 - 49579

  --1100000110101100    1100000110101101    1100000110101110    1100000110101111    1100000110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49580 - 49584

  --1100000110110001    1100000110110010    1100000110110011    1100000110110100    1100000110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49585 - 49589

  --1100000110110110    1100000110110111    1100000110111000    1100000110111001    1100000110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49590 - 49594

  --1100000110111011    1100000110111100    1100000110111101    1100000110111110    1100000110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49595 - 49599

  --1100000111000000    1100000111000001    1100000111000010    1100000111000011    1100000111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49600 - 49604

  --1100000111000101    1100000111000110    1100000111000111    1100000111001000    1100000111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49605 - 49609

  --1100000111001010    1100000111001011    1100000111001100    1100000111001101    1100000111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49610 - 49614

  --1100000111001111    1100000111010000    1100000111010001    1100000111010010    1100000111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49615 - 49619

  --1100000111010100    1100000111010101    1100000111010110    1100000111010111    1100000111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49620 - 49624

  --1100000111011001    1100000111011010    1100000111011011    1100000111011100    1100000111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49625 - 49629

  --1100000111011110    1100000111011111    1100000111100000    1100000111100001    1100000111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49630 - 49634

  --1100000111100011    1100000111100100    1100000111100101    1100000111100110    1100000111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49635 - 49639

  --1100000111101000    1100000111101001    1100000111101010    1100000111101011    1100000111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49640 - 49644

  --1100000111101101    1100000111101110    1100000111101111    1100000111110000    1100000111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49645 - 49649

  --1100000111110010    1100000111110011    1100000111110100    1100000111110101    1100000111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49650 - 49654

  --1100000111110111    1100000111111000    1100000111111001    1100000111111010    1100000111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49655 - 49659

  --1100000111111100    1100000111111101    1100000111111110    1100000111111111    1100001000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49660 - 49664

  --1100001000000001    1100001000000010    1100001000000011    1100001000000100    1100001000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49665 - 49669

  --1100001000000110    1100001000000111    1100001000001000    1100001000001001    1100001000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49670 - 49674

  --1100001000001011    1100001000001100    1100001000001101    1100001000001110    1100001000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49675 - 49679

  --1100001000010000    1100001000010001    1100001000010010    1100001000010011    1100001000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49680 - 49684

  --1100001000010101    1100001000010110    1100001000010111    1100001000011000    1100001000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49685 - 49689

  --1100001000011010    1100001000011011    1100001000011100    1100001000011101    1100001000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49690 - 49694

  --1100001000011111    1100001000100000    1100001000100001    1100001000100010    1100001000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49695 - 49699

  --1100001000100100    1100001000100101    1100001000100110    1100001000100111    1100001000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49700 - 49704

  --1100001000101001    1100001000101010    1100001000101011    1100001000101100    1100001000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49705 - 49709

  --1100001000101110    1100001000101111    1100001000110000    1100001000110001    1100001000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49710 - 49714

  --1100001000110011    1100001000110100    1100001000110101    1100001000110110    1100001000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49715 - 49719

  --1100001000111000    1100001000111001    1100001000111010    1100001000111011    1100001000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49720 - 49724

  --1100001000111101    1100001000111110    1100001000111111    1100001001000000    1100001001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49725 - 49729

  --1100001001000010    1100001001000011    1100001001000100    1100001001000101    1100001001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49730 - 49734

  --1100001001000111    1100001001001000    1100001001001001    1100001001001010    1100001001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49735 - 49739

  --1100001001001100    1100001001001101    1100001001001110    1100001001001111    1100001001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49740 - 49744

  --1100001001010001    1100001001010010    1100001001010011    1100001001010100    1100001001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49745 - 49749

  --1100001001010110    1100001001010111    1100001001011000    1100001001011001    1100001001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49750 - 49754

  --1100001001011011    1100001001011100    1100001001011101    1100001001011110    1100001001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49755 - 49759

  --1100001001100000    1100001001100001    1100001001100010    1100001001100011    1100001001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49760 - 49764

  --1100001001100101    1100001001100110    1100001001100111    1100001001101000    1100001001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49765 - 49769

  --1100001001101010    1100001001101011    1100001001101100    1100001001101101    1100001001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49770 - 49774

  --1100001001101111    1100001001110000    1100001001110001    1100001001110010    1100001001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49775 - 49779

  --1100001001110100    1100001001110101    1100001001110110    1100001001110111    1100001001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49780 - 49784

  --1100001001111001    1100001001111010    1100001001111011    1100001001111100    1100001001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49785 - 49789

  --1100001001111110    1100001001111111    1100001010000000    1100001010000001    1100001010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49790 - 49794

  --1100001010000011    1100001010000100    1100001010000101    1100001010000110    1100001010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49795 - 49799

  --1100001010001000    1100001010001001    1100001010001010    1100001010001011    1100001010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49800 - 49804

  --1100001010001101    1100001010001110    1100001010001111    1100001010010000    1100001010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49805 - 49809

  --1100001010010010    1100001010010011    1100001010010100    1100001010010101    1100001010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49810 - 49814

  --1100001010010111    1100001010011000    1100001010011001    1100001010011010    1100001010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49815 - 49819

  --1100001010011100    1100001010011101    1100001010011110    1100001010011111    1100001010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49820 - 49824

  --1100001010100001    1100001010100010    1100001010100011    1100001010100100    1100001010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49825 - 49829

  --1100001010100110    1100001010100111    1100001010101000    1100001010101001    1100001010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49830 - 49834

  --1100001010101011    1100001010101100    1100001010101101    1100001010101110    1100001010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49835 - 49839

  --1100001010110000    1100001010110001    1100001010110010    1100001010110011    1100001010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49840 - 49844

  --1100001010110101    1100001010110110    1100001010110111    1100001010111000    1100001010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49845 - 49849

  --1100001010111010    1100001010111011    1100001010111100    1100001010111101    1100001010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49850 - 49854

  --1100001010111111    1100001011000000    1100001011000001    1100001011000010    1100001011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49855 - 49859

  --1100001011000100    1100001011000101    1100001011000110    1100001011000111    1100001011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49860 - 49864

  --1100001011001001    1100001011001010    1100001011001011    1100001011001100    1100001011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49865 - 49869

  --1100001011001110    1100001011001111    1100001011010000    1100001011010001    1100001011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49870 - 49874

  --1100001011010011    1100001011010100    1100001011010101    1100001011010110    1100001011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49875 - 49879

  --1100001011011000    1100001011011001    1100001011011010    1100001011011011    1100001011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49880 - 49884

  --1100001011011101    1100001011011110    1100001011011111    1100001011100000    1100001011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49885 - 49889

  --1100001011100010    1100001011100011    1100001011100100    1100001011100101    1100001011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49890 - 49894

  --1100001011100111    1100001011101000    1100001011101001    1100001011101010    1100001011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49895 - 49899

  --1100001011101100    1100001011101101    1100001011101110    1100001011101111    1100001011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49900 - 49904

  --1100001011110001    1100001011110010    1100001011110011    1100001011110100    1100001011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49905 - 49909

  --1100001011110110    1100001011110111    1100001011111000    1100001011111001    1100001011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49910 - 49914

  --1100001011111011    1100001011111100    1100001011111101    1100001011111110    1100001011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49915 - 49919

  --1100001100000000    1100001100000001    1100001100000010    1100001100000011    1100001100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49920 - 49924

  --1100001100000101    1100001100000110    1100001100000111    1100001100001000    1100001100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49925 - 49929

  --1100001100001010    1100001100001011    1100001100001100    1100001100001101    1100001100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49930 - 49934

  --1100001100001111    1100001100010000    1100001100010001    1100001100010010    1100001100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49935 - 49939

  --1100001100010100    1100001100010101    1100001100010110    1100001100010111    1100001100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49940 - 49944

  --1100001100011001    1100001100011010    1100001100011011    1100001100011100    1100001100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49945 - 49949

  --1100001100011110    1100001100011111    1100001100100000    1100001100100001    1100001100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49950 - 49954

  --1100001100100011    1100001100100100    1100001100100101    1100001100100110    1100001100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49955 - 49959

  --1100001100101000    1100001100101001    1100001100101010    1100001100101011    1100001100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49960 - 49964

  --1100001100101101    1100001100101110    1100001100101111    1100001100110000    1100001100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49965 - 49969

  --1100001100110010    1100001100110011    1100001100110100    1100001100110101    1100001100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49970 - 49974

  --1100001100110111    1100001100111000    1100001100111001    1100001100111010    1100001100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49975 - 49979

  --1100001100111100    1100001100111101    1100001100111110    1100001100111111    1100001101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49980 - 49984

  --1100001101000001    1100001101000010    1100001101000011    1100001101000100    1100001101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49985 - 49989

  --1100001101000110    1100001101000111    1100001101001000    1100001101001001    1100001101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49990 - 49994

  --1100001101001011    1100001101001100    1100001101001101    1100001101001110    1100001101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 49995 - 49999

  --1100001101010000    1100001101010001    1100001101010010    1100001101010011    1100001101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50000 - 50004

  --1100001101010101    1100001101010110    1100001101010111    1100001101011000    1100001101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50005 - 50009

  --1100001101011010    1100001101011011    1100001101011100    1100001101011101    1100001101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50010 - 50014

  --1100001101011111    1100001101100000    1100001101100001    1100001101100010    1100001101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50015 - 50019

  --1100001101100100    1100001101100101    1100001101100110    1100001101100111    1100001101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50020 - 50024

  --1100001101101001    1100001101101010    1100001101101011    1100001101101100    1100001101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50025 - 50029

  --1100001101101110    1100001101101111    1100001101110000    1100001101110001    1100001101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50030 - 50034

  --1100001101110011    1100001101110100    1100001101110101    1100001101110110    1100001101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50035 - 50039

  --1100001101111000    1100001101111001    1100001101111010    1100001101111011    1100001101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50040 - 50044

  --1100001101111101    1100001101111110    1100001101111111    1100001110000000    1100001110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50045 - 50049

  --1100001110000010    1100001110000011    1100001110000100    1100001110000101    1100001110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50050 - 50054

  --1100001110000111    1100001110001000    1100001110001001    1100001110001010    1100001110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50055 - 50059

  --1100001110001100    1100001110001101    1100001110001110    1100001110001111    1100001110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50060 - 50064

  --1100001110010001    1100001110010010    1100001110010011    1100001110010100    1100001110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50065 - 50069

  --1100001110010110    1100001110010111    1100001110011000    1100001110011001    1100001110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50070 - 50074

  --1100001110011011    1100001110011100    1100001110011101    1100001110011110    1100001110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50075 - 50079

  --1100001110100000    1100001110100001    1100001110100010    1100001110100011    1100001110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50080 - 50084

  --1100001110100101    1100001110100110    1100001110100111    1100001110101000    1100001110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50085 - 50089

  --1100001110101010    1100001110101011    1100001110101100    1100001110101101    1100001110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50090 - 50094

  --1100001110101111    1100001110110000    1100001110110001    1100001110110010    1100001110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50095 - 50099

  --1100001110110100    1100001110110101    1100001110110110    1100001110110111    1100001110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50100 - 50104

  --1100001110111001    1100001110111010    1100001110111011    1100001110111100    1100001110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50105 - 50109

  --1100001110111110    1100001110111111    1100001111000000    1100001111000001    1100001111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50110 - 50114

  --1100001111000011    1100001111000100    1100001111000101    1100001111000110    1100001111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50115 - 50119

  --1100001111001000    1100001111001001    1100001111001010    1100001111001011    1100001111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50120 - 50124

  --1100001111001101    1100001111001110    1100001111001111    1100001111010000    1100001111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50125 - 50129

  --1100001111010010    1100001111010011    1100001111010100    1100001111010101    1100001111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50130 - 50134

  --1100001111010111    1100001111011000    1100001111011001    1100001111011010    1100001111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50135 - 50139

  --1100001111011100    1100001111011101    1100001111011110    1100001111011111    1100001111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50140 - 50144

  --1100001111100001    1100001111100010    1100001111100011    1100001111100100    1100001111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50145 - 50149

  --1100001111100110    1100001111100111    1100001111101000    1100001111101001    1100001111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50150 - 50154

  --1100001111101011    1100001111101100    1100001111101101    1100001111101110    1100001111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50155 - 50159

  --1100001111110000    1100001111110001    1100001111110010    1100001111110011    1100001111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50160 - 50164

  --1100001111110101    1100001111110110    1100001111110111    1100001111111000    1100001111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50165 - 50169

  --1100001111111010    1100001111111011    1100001111111100    1100001111111101    1100001111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50170 - 50174

  --1100001111111111    1100010000000000    1100010000000001    1100010000000010    1100010000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50175 - 50179

  --1100010000000100    1100010000000101    1100010000000110    1100010000000111    1100010000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50180 - 50184

  --1100010000001001    1100010000001010    1100010000001011    1100010000001100    1100010000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50185 - 50189

  --1100010000001110    1100010000001111    1100010000010000    1100010000010001    1100010000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50190 - 50194

  --1100010000010011    1100010000010100    1100010000010101    1100010000010110    1100010000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50195 - 50199

  --1100010000011000    1100010000011001    1100010000011010    1100010000011011    1100010000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50200 - 50204

  --1100010000011101    1100010000011110    1100010000011111    1100010000100000    1100010000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50205 - 50209

  --1100010000100010    1100010000100011    1100010000100100    1100010000100101    1100010000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50210 - 50214

  --1100010000100111    1100010000101000    1100010000101001    1100010000101010    1100010000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50215 - 50219

  --1100010000101100    1100010000101101    1100010000101110    1100010000101111    1100010000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50220 - 50224

  --1100010000110001    1100010000110010    1100010000110011    1100010000110100    1100010000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50225 - 50229

  --1100010000110110    1100010000110111    1100010000111000    1100010000111001    1100010000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50230 - 50234

  --1100010000111011    1100010000111100    1100010000111101    1100010000111110    1100010000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50235 - 50239

  --1100010001000000    1100010001000001    1100010001000010    1100010001000011    1100010001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50240 - 50244

  --1100010001000101    1100010001000110    1100010001000111    1100010001001000    1100010001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50245 - 50249

  --1100010001001010    1100010001001011    1100010001001100    1100010001001101    1100010001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50250 - 50254

  --1100010001001111    1100010001010000    1100010001010001    1100010001010010    1100010001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50255 - 50259

  --1100010001010100    1100010001010101    1100010001010110    1100010001010111    1100010001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50260 - 50264

  --1100010001011001    1100010001011010    1100010001011011    1100010001011100    1100010001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50265 - 50269

  --1100010001011110    1100010001011111    1100010001100000    1100010001100001    1100010001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50270 - 50274

  --1100010001100011    1100010001100100    1100010001100101    1100010001100110    1100010001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50275 - 50279

  --1100010001101000    1100010001101001    1100010001101010    1100010001101011    1100010001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50280 - 50284

  --1100010001101101    1100010001101110    1100010001101111    1100010001110000    1100010001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50285 - 50289

  --1100010001110010    1100010001110011    1100010001110100    1100010001110101    1100010001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50290 - 50294

  --1100010001110111    1100010001111000    1100010001111001    1100010001111010    1100010001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50295 - 50299

  --1100010001111100    1100010001111101    1100010001111110    1100010001111111    1100010010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50300 - 50304

  --1100010010000001    1100010010000010    1100010010000011    1100010010000100    1100010010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50305 - 50309

  --1100010010000110    1100010010000111    1100010010001000    1100010010001001    1100010010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50310 - 50314

  --1100010010001011    1100010010001100    1100010010001101    1100010010001110    1100010010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50315 - 50319

  --1100010010010000    1100010010010001    1100010010010010    1100010010010011    1100010010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50320 - 50324

  --1100010010010101    1100010010010110    1100010010010111    1100010010011000    1100010010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50325 - 50329

  --1100010010011010    1100010010011011    1100010010011100    1100010010011101    1100010010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50330 - 50334

  --1100010010011111    1100010010100000    1100010010100001    1100010010100010    1100010010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50335 - 50339

  --1100010010100100    1100010010100101    1100010010100110    1100010010100111    1100010010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50340 - 50344

  --1100010010101001    1100010010101010    1100010010101011    1100010010101100    1100010010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50345 - 50349

  --1100010010101110    1100010010101111    1100010010110000    1100010010110001    1100010010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50350 - 50354

  --1100010010110011    1100010010110100    1100010010110101    1100010010110110    1100010010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50355 - 50359

  --1100010010111000    1100010010111001    1100010010111010    1100010010111011    1100010010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50360 - 50364

  --1100010010111101    1100010010111110    1100010010111111    1100010011000000    1100010011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50365 - 50369

  --1100010011000010    1100010011000011    1100010011000100    1100010011000101    1100010011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50370 - 50374

  --1100010011000111    1100010011001000    1100010011001001    1100010011001010    1100010011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50375 - 50379

  --1100010011001100    1100010011001101    1100010011001110    1100010011001111    1100010011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50380 - 50384

  --1100010011010001    1100010011010010    1100010011010011    1100010011010100    1100010011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50385 - 50389

  --1100010011010110    1100010011010111    1100010011011000    1100010011011001    1100010011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50390 - 50394

  --1100010011011011    1100010011011100    1100010011011101    1100010011011110    1100010011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50395 - 50399

  --1100010011100000    1100010011100001    1100010011100010    1100010011100011    1100010011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50400 - 50404

  --1100010011100101    1100010011100110    1100010011100111    1100010011101000    1100010011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50405 - 50409

  --1100010011101010    1100010011101011    1100010011101100    1100010011101101    1100010011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50410 - 50414

  --1100010011101111    1100010011110000    1100010011110001    1100010011110010    1100010011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50415 - 50419

  --1100010011110100    1100010011110101    1100010011110110    1100010011110111    1100010011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50420 - 50424

  --1100010011111001    1100010011111010    1100010011111011    1100010011111100    1100010011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50425 - 50429

  --1100010011111110    1100010011111111    1100010100000000    1100010100000001    1100010100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50430 - 50434

  --1100010100000011    1100010100000100    1100010100000101    1100010100000110    1100010100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50435 - 50439

  --1100010100001000    1100010100001001    1100010100001010    1100010100001011    1100010100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50440 - 50444

  --1100010100001101    1100010100001110    1100010100001111    1100010100010000    1100010100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50445 - 50449

  --1100010100010010    1100010100010011    1100010100010100    1100010100010101    1100010100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50450 - 50454

  --1100010100010111    1100010100011000    1100010100011001    1100010100011010    1100010100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50455 - 50459

  --1100010100011100    1100010100011101    1100010100011110    1100010100011111    1100010100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50460 - 50464

  --1100010100100001    1100010100100010    1100010100100011    1100010100100100    1100010100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50465 - 50469

  --1100010100100110    1100010100100111    1100010100101000    1100010100101001    1100010100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50470 - 50474

  --1100010100101011    1100010100101100    1100010100101101    1100010100101110    1100010100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50475 - 50479

  --1100010100110000    1100010100110001    1100010100110010    1100010100110011    1100010100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50480 - 50484

  --1100010100110101    1100010100110110    1100010100110111    1100010100111000    1100010100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50485 - 50489

  --1100010100111010    1100010100111011    1100010100111100    1100010100111101    1100010100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50490 - 50494

  --1100010100111111    1100010101000000    1100010101000001    1100010101000010    1100010101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50495 - 50499

  --1100010101000100    1100010101000101    1100010101000110    1100010101000111    1100010101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50500 - 50504

  --1100010101001001    1100010101001010    1100010101001011    1100010101001100    1100010101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50505 - 50509

  --1100010101001110    1100010101001111    1100010101010000    1100010101010001    1100010101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50510 - 50514

  --1100010101010011    1100010101010100    1100010101010101    1100010101010110    1100010101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50515 - 50519

  --1100010101011000    1100010101011001    1100010101011010    1100010101011011    1100010101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50520 - 50524

  --1100010101011101    1100010101011110    1100010101011111    1100010101100000    1100010101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50525 - 50529

  --1100010101100010    1100010101100011    1100010101100100    1100010101100101    1100010101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50530 - 50534

  --1100010101100111    1100010101101000    1100010101101001    1100010101101010    1100010101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50535 - 50539

  --1100010101101100    1100010101101101    1100010101101110    1100010101101111    1100010101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50540 - 50544

  --1100010101110001    1100010101110010    1100010101110011    1100010101110100    1100010101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50545 - 50549

  --1100010101110110    1100010101110111    1100010101111000    1100010101111001    1100010101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50550 - 50554

  --1100010101111011    1100010101111100    1100010101111101    1100010101111110    1100010101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50555 - 50559

  --1100010110000000    1100010110000001    1100010110000010    1100010110000011    1100010110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50560 - 50564

  --1100010110000101    1100010110000110    1100010110000111    1100010110001000    1100010110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50565 - 50569

  --1100010110001010    1100010110001011    1100010110001100    1100010110001101    1100010110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50570 - 50574

  --1100010110001111    1100010110010000    1100010110010001    1100010110010010    1100010110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50575 - 50579

  --1100010110010100    1100010110010101    1100010110010110    1100010110010111    1100010110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50580 - 50584

  --1100010110011001    1100010110011010    1100010110011011    1100010110011100    1100010110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50585 - 50589

  --1100010110011110    1100010110011111    1100010110100000    1100010110100001    1100010110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50590 - 50594

  --1100010110100011    1100010110100100    1100010110100101    1100010110100110    1100010110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50595 - 50599

  --1100010110101000    1100010110101001    1100010110101010    1100010110101011    1100010110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50600 - 50604

  --1100010110101101    1100010110101110    1100010110101111    1100010110110000    1100010110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50605 - 50609

  --1100010110110010    1100010110110011    1100010110110100    1100010110110101    1100010110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50610 - 50614

  --1100010110110111    1100010110111000    1100010110111001    1100010110111010    1100010110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50615 - 50619

  --1100010110111100    1100010110111101    1100010110111110    1100010110111111    1100010111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50620 - 50624

  --1100010111000001    1100010111000010    1100010111000011    1100010111000100    1100010111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50625 - 50629

  --1100010111000110    1100010111000111    1100010111001000    1100010111001001    1100010111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50630 - 50634

  --1100010111001011    1100010111001100    1100010111001101    1100010111001110    1100010111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50635 - 50639

  --1100010111010000    1100010111010001    1100010111010010    1100010111010011    1100010111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50640 - 50644

  --1100010111010101    1100010111010110    1100010111010111    1100010111011000    1100010111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50645 - 50649

  --1100010111011010    1100010111011011    1100010111011100    1100010111011101    1100010111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50650 - 50654

  --1100010111011111    1100010111100000    1100010111100001    1100010111100010    1100010111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50655 - 50659

  --1100010111100100    1100010111100101    1100010111100110    1100010111100111    1100010111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50660 - 50664

  --1100010111101001    1100010111101010    1100010111101011    1100010111101100    1100010111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50665 - 50669

  --1100010111101110    1100010111101111    1100010111110000    1100010111110001    1100010111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50670 - 50674

  --1100010111110011    1100010111110100    1100010111110101    1100010111110110    1100010111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50675 - 50679

  --1100010111111000    1100010111111001    1100010111111010    1100010111111011    1100010111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50680 - 50684

  --1100010111111101    1100010111111110    1100010111111111    1100011000000000    1100011000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50685 - 50689

  --1100011000000010    1100011000000011    1100011000000100    1100011000000101    1100011000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50690 - 50694

  --1100011000000111    1100011000001000    1100011000001001    1100011000001010    1100011000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50695 - 50699

  --1100011000001100    1100011000001101    1100011000001110    1100011000001111    1100011000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50700 - 50704

  --1100011000010001    1100011000010010    1100011000010011    1100011000010100    1100011000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50705 - 50709

  --1100011000010110    1100011000010111    1100011000011000    1100011000011001    1100011000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50710 - 50714

  --1100011000011011    1100011000011100    1100011000011101    1100011000011110    1100011000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50715 - 50719

  --1100011000100000    1100011000100001    1100011000100010    1100011000100011    1100011000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50720 - 50724

  --1100011000100101    1100011000100110    1100011000100111    1100011000101000    1100011000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50725 - 50729

  --1100011000101010    1100011000101011    1100011000101100    1100011000101101    1100011000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50730 - 50734

  --1100011000101111    1100011000110000    1100011000110001    1100011000110010    1100011000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50735 - 50739

  --1100011000110100    1100011000110101    1100011000110110    1100011000110111    1100011000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50740 - 50744

  --1100011000111001    1100011000111010    1100011000111011    1100011000111100    1100011000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50745 - 50749

  --1100011000111110    1100011000111111    1100011001000000    1100011001000001    1100011001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50750 - 50754

  --1100011001000011    1100011001000100    1100011001000101    1100011001000110    1100011001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50755 - 50759

  --1100011001001000    1100011001001001    1100011001001010    1100011001001011    1100011001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50760 - 50764

  --1100011001001101    1100011001001110    1100011001001111    1100011001010000    1100011001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50765 - 50769

  --1100011001010010    1100011001010011    1100011001010100    1100011001010101    1100011001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50770 - 50774

  --1100011001010111    1100011001011000    1100011001011001    1100011001011010    1100011001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50775 - 50779

  --1100011001011100    1100011001011101    1100011001011110    1100011001011111    1100011001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50780 - 50784

  --1100011001100001    1100011001100010    1100011001100011    1100011001100100    1100011001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50785 - 50789

  --1100011001100110    1100011001100111    1100011001101000    1100011001101001    1100011001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50790 - 50794

  --1100011001101011    1100011001101100    1100011001101101    1100011001101110    1100011001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50795 - 50799

  --1100011001110000    1100011001110001    1100011001110010    1100011001110011    1100011001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50800 - 50804

  --1100011001110101    1100011001110110    1100011001110111    1100011001111000    1100011001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50805 - 50809

  --1100011001111010    1100011001111011    1100011001111100    1100011001111101    1100011001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50810 - 50814

  --1100011001111111    1100011010000000    1100011010000001    1100011010000010    1100011010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50815 - 50819

  --1100011010000100    1100011010000101    1100011010000110    1100011010000111    1100011010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50820 - 50824

  --1100011010001001    1100011010001010    1100011010001011    1100011010001100    1100011010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50825 - 50829

  --1100011010001110    1100011010001111    1100011010010000    1100011010010001    1100011010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50830 - 50834

  --1100011010010011    1100011010010100    1100011010010101    1100011010010110    1100011010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50835 - 50839

  --1100011010011000    1100011010011001    1100011010011010    1100011010011011    1100011010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50840 - 50844

  --1100011010011101    1100011010011110    1100011010011111    1100011010100000    1100011010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50845 - 50849

  --1100011010100010    1100011010100011    1100011010100100    1100011010100101    1100011010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50850 - 50854

  --1100011010100111    1100011010101000    1100011010101001    1100011010101010    1100011010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50855 - 50859

  --1100011010101100    1100011010101101    1100011010101110    1100011010101111    1100011010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50860 - 50864

  --1100011010110001    1100011010110010    1100011010110011    1100011010110100    1100011010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50865 - 50869

  --1100011010110110    1100011010110111    1100011010111000    1100011010111001    1100011010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50870 - 50874

  --1100011010111011    1100011010111100    1100011010111101    1100011010111110    1100011010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50875 - 50879

  --1100011011000000    1100011011000001    1100011011000010    1100011011000011    1100011011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50880 - 50884

  --1100011011000101    1100011011000110    1100011011000111    1100011011001000    1100011011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50885 - 50889

  --1100011011001010    1100011011001011    1100011011001100    1100011011001101    1100011011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50890 - 50894

  --1100011011001111    1100011011010000    1100011011010001    1100011011010010    1100011011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50895 - 50899

  --1100011011010100    1100011011010101    1100011011010110    1100011011010111    1100011011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50900 - 50904

  --1100011011011001    1100011011011010    1100011011011011    1100011011011100    1100011011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50905 - 50909

  --1100011011011110    1100011011011111    1100011011100000    1100011011100001    1100011011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50910 - 50914

  --1100011011100011    1100011011100100    1100011011100101    1100011011100110    1100011011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50915 - 50919

  --1100011011101000    1100011011101001    1100011011101010    1100011011101011    1100011011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50920 - 50924

  --1100011011101101    1100011011101110    1100011011101111    1100011011110000    1100011011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50925 - 50929

  --1100011011110010    1100011011110011    1100011011110100    1100011011110101    1100011011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50930 - 50934

  --1100011011110111    1100011011111000    1100011011111001    1100011011111010    1100011011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50935 - 50939

  --1100011011111100    1100011011111101    1100011011111110    1100011011111111    1100011100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50940 - 50944

  --1100011100000001    1100011100000010    1100011100000011    1100011100000100    1100011100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50945 - 50949

  --1100011100000110    1100011100000111    1100011100001000    1100011100001001    1100011100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50950 - 50954

  --1100011100001011    1100011100001100    1100011100001101    1100011100001110    1100011100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50955 - 50959

  --1100011100010000    1100011100010001    1100011100010010    1100011100010011    1100011100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50960 - 50964

  --1100011100010101    1100011100010110    1100011100010111    1100011100011000    1100011100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50965 - 50969

  --1100011100011010    1100011100011011    1100011100011100    1100011100011101    1100011100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50970 - 50974

  --1100011100011111    1100011100100000    1100011100100001    1100011100100010    1100011100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50975 - 50979

  --1100011100100100    1100011100100101    1100011100100110    1100011100100111    1100011100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50980 - 50984

  --1100011100101001    1100011100101010    1100011100101011    1100011100101100    1100011100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50985 - 50989

  --1100011100101110    1100011100101111    1100011100110000    1100011100110001    1100011100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50990 - 50994

  --1100011100110011    1100011100110100    1100011100110101    1100011100110110    1100011100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 50995 - 50999

  --1100011100111000    1100011100111001    1100011100111010    1100011100111011    1100011100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51000 - 51004

  --1100011100111101    1100011100111110    1100011100111111    1100011101000000    1100011101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51005 - 51009

  --1100011101000010    1100011101000011    1100011101000100    1100011101000101    1100011101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51010 - 51014

  --1100011101000111    1100011101001000    1100011101001001    1100011101001010    1100011101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51015 - 51019

  --1100011101001100    1100011101001101    1100011101001110    1100011101001111    1100011101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51020 - 51024

  --1100011101010001    1100011101010010    1100011101010011    1100011101010100    1100011101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51025 - 51029

  --1100011101010110    1100011101010111    1100011101011000    1100011101011001    1100011101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51030 - 51034

  --1100011101011011    1100011101011100    1100011101011101    1100011101011110    1100011101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51035 - 51039

  --1100011101100000    1100011101100001    1100011101100010    1100011101100011    1100011101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51040 - 51044

  --1100011101100101    1100011101100110    1100011101100111    1100011101101000    1100011101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51045 - 51049

  --1100011101101010    1100011101101011    1100011101101100    1100011101101101    1100011101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51050 - 51054

  --1100011101101111    1100011101110000    1100011101110001    1100011101110010    1100011101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51055 - 51059

  --1100011101110100    1100011101110101    1100011101110110    1100011101110111    1100011101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51060 - 51064

  --1100011101111001    1100011101111010    1100011101111011    1100011101111100    1100011101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51065 - 51069

  --1100011101111110    1100011101111111    1100011110000000    1100011110000001    1100011110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51070 - 51074

  --1100011110000011    1100011110000100    1100011110000101    1100011110000110    1100011110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51075 - 51079

  --1100011110001000    1100011110001001    1100011110001010    1100011110001011    1100011110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51080 - 51084

  --1100011110001101    1100011110001110    1100011110001111    1100011110010000    1100011110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51085 - 51089

  --1100011110010010    1100011110010011    1100011110010100    1100011110010101    1100011110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51090 - 51094

  --1100011110010111    1100011110011000    1100011110011001    1100011110011010    1100011110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51095 - 51099

  --1100011110011100    1100011110011101    1100011110011110    1100011110011111    1100011110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51100 - 51104

  --1100011110100001    1100011110100010    1100011110100011    1100011110100100    1100011110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51105 - 51109

  --1100011110100110    1100011110100111    1100011110101000    1100011110101001    1100011110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51110 - 51114

  --1100011110101011    1100011110101100    1100011110101101    1100011110101110    1100011110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51115 - 51119

  --1100011110110000    1100011110110001    1100011110110010    1100011110110011    1100011110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51120 - 51124

  --1100011110110101    1100011110110110    1100011110110111    1100011110111000    1100011110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51125 - 51129

  --1100011110111010    1100011110111011    1100011110111100    1100011110111101    1100011110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51130 - 51134

  --1100011110111111    1100011111000000    1100011111000001    1100011111000010    1100011111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51135 - 51139

  --1100011111000100    1100011111000101    1100011111000110    1100011111000111    1100011111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51140 - 51144

  --1100011111001001    1100011111001010    1100011111001011    1100011111001100    1100011111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51145 - 51149

  --1100011111001110    1100011111001111    1100011111010000    1100011111010001    1100011111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51150 - 51154

  --1100011111010011    1100011111010100    1100011111010101    1100011111010110    1100011111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51155 - 51159

  --1100011111011000    1100011111011001    1100011111011010    1100011111011011    1100011111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51160 - 51164

  --1100011111011101    1100011111011110    1100011111011111    1100011111100000    1100011111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51165 - 51169

  --1100011111100010    1100011111100011    1100011111100100    1100011111100101    1100011111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51170 - 51174

  --1100011111100111    1100011111101000    1100011111101001    1100011111101010    1100011111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51175 - 51179

  --1100011111101100    1100011111101101    1100011111101110    1100011111101111    1100011111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51180 - 51184

  --1100011111110001    1100011111110010    1100011111110011    1100011111110100    1100011111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51185 - 51189

  --1100011111110110    1100011111110111    1100011111111000    1100011111111001    1100011111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51190 - 51194

  --1100011111111011    1100011111111100    1100011111111101    1100011111111110    1100011111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51195 - 51199

  --1100100000000000    1100100000000001    1100100000000010    1100100000000011    1100100000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51200 - 51204

  --1100100000000101    1100100000000110    1100100000000111    1100100000001000    1100100000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51205 - 51209

  --1100100000001010    1100100000001011    1100100000001100    1100100000001101    1100100000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51210 - 51214

  --1100100000001111    1100100000010000    1100100000010001    1100100000010010    1100100000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51215 - 51219

  --1100100000010100    1100100000010101    1100100000010110    1100100000010111    1100100000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51220 - 51224

  --1100100000011001    1100100000011010    1100100000011011    1100100000011100    1100100000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51225 - 51229

  --1100100000011110    1100100000011111    1100100000100000    1100100000100001    1100100000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51230 - 51234

  --1100100000100011    1100100000100100    1100100000100101    1100100000100110    1100100000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51235 - 51239

  --1100100000101000    1100100000101001    1100100000101010    1100100000101011    1100100000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51240 - 51244

  --1100100000101101    1100100000101110    1100100000101111    1100100000110000    1100100000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51245 - 51249

  --1100100000110010    1100100000110011    1100100000110100    1100100000110101    1100100000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51250 - 51254

  --1100100000110111    1100100000111000    1100100000111001    1100100000111010    1100100000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51255 - 51259

  --1100100000111100    1100100000111101    1100100000111110    1100100000111111    1100100001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51260 - 51264

  --1100100001000001    1100100001000010    1100100001000011    1100100001000100    1100100001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51265 - 51269

  --1100100001000110    1100100001000111    1100100001001000    1100100001001001    1100100001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51270 - 51274

  --1100100001001011    1100100001001100    1100100001001101    1100100001001110    1100100001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51275 - 51279

  --1100100001010000    1100100001010001    1100100001010010    1100100001010011    1100100001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51280 - 51284

  --1100100001010101    1100100001010110    1100100001010111    1100100001011000    1100100001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51285 - 51289

  --1100100001011010    1100100001011011    1100100001011100    1100100001011101    1100100001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51290 - 51294

  --1100100001011111    1100100001100000    1100100001100001    1100100001100010    1100100001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51295 - 51299

  --1100100001100100    1100100001100101    1100100001100110    1100100001100111    1100100001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51300 - 51304

  --1100100001101001    1100100001101010    1100100001101011    1100100001101100    1100100001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51305 - 51309

  --1100100001101110    1100100001101111    1100100001110000    1100100001110001    1100100001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51310 - 51314

  --1100100001110011    1100100001110100    1100100001110101    1100100001110110    1100100001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51315 - 51319

  --1100100001111000    1100100001111001    1100100001111010    1100100001111011    1100100001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51320 - 51324

  --1100100001111101    1100100001111110    1100100001111111    1100100010000000    1100100010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51325 - 51329

  --1100100010000010    1100100010000011    1100100010000100    1100100010000101    1100100010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51330 - 51334

  --1100100010000111    1100100010001000    1100100010001001    1100100010001010    1100100010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51335 - 51339

  --1100100010001100    1100100010001101    1100100010001110    1100100010001111    1100100010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51340 - 51344

  --1100100010010001    1100100010010010    1100100010010011    1100100010010100    1100100010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51345 - 51349

  --1100100010010110    1100100010010111    1100100010011000    1100100010011001    1100100010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51350 - 51354

  --1100100010011011    1100100010011100    1100100010011101    1100100010011110    1100100010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51355 - 51359

  --1100100010100000    1100100010100001    1100100010100010    1100100010100011    1100100010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51360 - 51364

  --1100100010100101    1100100010100110    1100100010100111    1100100010101000    1100100010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51365 - 51369

  --1100100010101010    1100100010101011    1100100010101100    1100100010101101    1100100010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51370 - 51374

  --1100100010101111    1100100010110000    1100100010110001    1100100010110010    1100100010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51375 - 51379

  --1100100010110100    1100100010110101    1100100010110110    1100100010110111    1100100010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51380 - 51384

  --1100100010111001    1100100010111010    1100100010111011    1100100010111100    1100100010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51385 - 51389

  --1100100010111110    1100100010111111    1100100011000000    1100100011000001    1100100011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51390 - 51394

  --1100100011000011    1100100011000100    1100100011000101    1100100011000110    1100100011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51395 - 51399

  --1100100011001000    1100100011001001    1100100011001010    1100100011001011    1100100011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51400 - 51404

  --1100100011001101    1100100011001110    1100100011001111    1100100011010000    1100100011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51405 - 51409

  --1100100011010010    1100100011010011    1100100011010100    1100100011010101    1100100011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51410 - 51414

  --1100100011010111    1100100011011000    1100100011011001    1100100011011010    1100100011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51415 - 51419

  --1100100011011100    1100100011011101    1100100011011110    1100100011011111    1100100011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51420 - 51424

  --1100100011100001    1100100011100010    1100100011100011    1100100011100100    1100100011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51425 - 51429

  --1100100011100110    1100100011100111    1100100011101000    1100100011101001    1100100011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51430 - 51434

  --1100100011101011    1100100011101100    1100100011101101    1100100011101110    1100100011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51435 - 51439

  --1100100011110000    1100100011110001    1100100011110010    1100100011110011    1100100011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51440 - 51444

  --1100100011110101    1100100011110110    1100100011110111    1100100011111000    1100100011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51445 - 51449

  --1100100011111010    1100100011111011    1100100011111100    1100100011111101    1100100011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51450 - 51454

  --1100100011111111    1100100100000000    1100100100000001    1100100100000010    1100100100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51455 - 51459

  --1100100100000100    1100100100000101    1100100100000110    1100100100000111    1100100100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51460 - 51464

  --1100100100001001    1100100100001010    1100100100001011    1100100100001100    1100100100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51465 - 51469

  --1100100100001110    1100100100001111    1100100100010000    1100100100010001    1100100100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51470 - 51474

  --1100100100010011    1100100100010100    1100100100010101    1100100100010110    1100100100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51475 - 51479

  --1100100100011000    1100100100011001    1100100100011010    1100100100011011    1100100100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51480 - 51484

  --1100100100011101    1100100100011110    1100100100011111    1100100100100000    1100100100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51485 - 51489

  --1100100100100010    1100100100100011    1100100100100100    1100100100100101    1100100100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51490 - 51494

  --1100100100100111    1100100100101000    1100100100101001    1100100100101010    1100100100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51495 - 51499

  --1100100100101100    1100100100101101    1100100100101110    1100100100101111    1100100100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51500 - 51504

  --1100100100110001    1100100100110010    1100100100110011    1100100100110100    1100100100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51505 - 51509

  --1100100100110110    1100100100110111    1100100100111000    1100100100111001    1100100100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51510 - 51514

  --1100100100111011    1100100100111100    1100100100111101    1100100100111110    1100100100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51515 - 51519

  --1100100101000000    1100100101000001    1100100101000010    1100100101000011    1100100101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51520 - 51524

  --1100100101000101    1100100101000110    1100100101000111    1100100101001000    1100100101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51525 - 51529

  --1100100101001010    1100100101001011    1100100101001100    1100100101001101    1100100101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51530 - 51534

  --1100100101001111    1100100101010000    1100100101010001    1100100101010010    1100100101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51535 - 51539

  --1100100101010100    1100100101010101    1100100101010110    1100100101010111    1100100101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51540 - 51544

  --1100100101011001    1100100101011010    1100100101011011    1100100101011100    1100100101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51545 - 51549

  --1100100101011110    1100100101011111    1100100101100000    1100100101100001    1100100101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51550 - 51554

  --1100100101100011    1100100101100100    1100100101100101    1100100101100110    1100100101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51555 - 51559

  --1100100101101000    1100100101101001    1100100101101010    1100100101101011    1100100101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51560 - 51564

  --1100100101101101    1100100101101110    1100100101101111    1100100101110000    1100100101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51565 - 51569

  --1100100101110010    1100100101110011    1100100101110100    1100100101110101    1100100101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51570 - 51574

  --1100100101110111    1100100101111000    1100100101111001    1100100101111010    1100100101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51575 - 51579

  --1100100101111100    1100100101111101    1100100101111110    1100100101111111    1100100110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51580 - 51584

  --1100100110000001    1100100110000010    1100100110000011    1100100110000100    1100100110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51585 - 51589

  --1100100110000110    1100100110000111    1100100110001000    1100100110001001    1100100110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51590 - 51594

  --1100100110001011    1100100110001100    1100100110001101    1100100110001110    1100100110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51595 - 51599

  --1100100110010000    1100100110010001    1100100110010010    1100100110010011    1100100110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51600 - 51604

  --1100100110010101    1100100110010110    1100100110010111    1100100110011000    1100100110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51605 - 51609

  --1100100110011010    1100100110011011    1100100110011100    1100100110011101    1100100110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51610 - 51614

  --1100100110011111    1100100110100000    1100100110100001    1100100110100010    1100100110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51615 - 51619

  --1100100110100100    1100100110100101    1100100110100110    1100100110100111    1100100110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51620 - 51624

  --1100100110101001    1100100110101010    1100100110101011    1100100110101100    1100100110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51625 - 51629

  --1100100110101110    1100100110101111    1100100110110000    1100100110110001    1100100110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51630 - 51634

  --1100100110110011    1100100110110100    1100100110110101    1100100110110110    1100100110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51635 - 51639

  --1100100110111000    1100100110111001    1100100110111010    1100100110111011    1100100110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51640 - 51644

  --1100100110111101    1100100110111110    1100100110111111    1100100111000000    1100100111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51645 - 51649

  --1100100111000010    1100100111000011    1100100111000100    1100100111000101    1100100111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51650 - 51654

  --1100100111000111    1100100111001000    1100100111001001    1100100111001010    1100100111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51655 - 51659

  --1100100111001100    1100100111001101    1100100111001110    1100100111001111    1100100111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51660 - 51664

  --1100100111010001    1100100111010010    1100100111010011    1100100111010100    1100100111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51665 - 51669

  --1100100111010110    1100100111010111    1100100111011000    1100100111011001    1100100111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51670 - 51674

  --1100100111011011    1100100111011100    1100100111011101    1100100111011110    1100100111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51675 - 51679

  --1100100111100000    1100100111100001    1100100111100010    1100100111100011    1100100111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51680 - 51684

  --1100100111100101    1100100111100110    1100100111100111    1100100111101000    1100100111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51685 - 51689

  --1100100111101010    1100100111101011    1100100111101100    1100100111101101    1100100111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51690 - 51694

  --1100100111101111    1100100111110000    1100100111110001    1100100111110010    1100100111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51695 - 51699

  --1100100111110100    1100100111110101    1100100111110110    1100100111110111    1100100111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51700 - 51704

  --1100100111111001    1100100111111010    1100100111111011    1100100111111100    1100100111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51705 - 51709

  --1100100111111110    1100100111111111    1100101000000000    1100101000000001    1100101000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51710 - 51714

  --1100101000000011    1100101000000100    1100101000000101    1100101000000110    1100101000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51715 - 51719

  --1100101000001000    1100101000001001    1100101000001010    1100101000001011    1100101000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51720 - 51724

  --1100101000001101    1100101000001110    1100101000001111    1100101000010000    1100101000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51725 - 51729

  --1100101000010010    1100101000010011    1100101000010100    1100101000010101    1100101000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51730 - 51734

  --1100101000010111    1100101000011000    1100101000011001    1100101000011010    1100101000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51735 - 51739

  --1100101000011100    1100101000011101    1100101000011110    1100101000011111    1100101000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51740 - 51744

  --1100101000100001    1100101000100010    1100101000100011    1100101000100100    1100101000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51745 - 51749

  --1100101000100110    1100101000100111    1100101000101000    1100101000101001    1100101000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51750 - 51754

  --1100101000101011    1100101000101100    1100101000101101    1100101000101110    1100101000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51755 - 51759

  --1100101000110000    1100101000110001    1100101000110010    1100101000110011    1100101000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51760 - 51764

  --1100101000110101    1100101000110110    1100101000110111    1100101000111000    1100101000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51765 - 51769

  --1100101000111010    1100101000111011    1100101000111100    1100101000111101    1100101000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51770 - 51774

  --1100101000111111    1100101001000000    1100101001000001    1100101001000010    1100101001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51775 - 51779

  --1100101001000100    1100101001000101    1100101001000110    1100101001000111    1100101001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51780 - 51784

  --1100101001001001    1100101001001010    1100101001001011    1100101001001100    1100101001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51785 - 51789

  --1100101001001110    1100101001001111    1100101001010000    1100101001010001    1100101001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51790 - 51794

  --1100101001010011    1100101001010100    1100101001010101    1100101001010110    1100101001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51795 - 51799

  --1100101001011000    1100101001011001    1100101001011010    1100101001011011    1100101001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51800 - 51804

  --1100101001011101    1100101001011110    1100101001011111    1100101001100000    1100101001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51805 - 51809

  --1100101001100010    1100101001100011    1100101001100100    1100101001100101    1100101001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51810 - 51814

  --1100101001100111    1100101001101000    1100101001101001    1100101001101010    1100101001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51815 - 51819

  --1100101001101100    1100101001101101    1100101001101110    1100101001101111    1100101001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51820 - 51824

  --1100101001110001    1100101001110010    1100101001110011    1100101001110100    1100101001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51825 - 51829

  --1100101001110110    1100101001110111    1100101001111000    1100101001111001    1100101001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51830 - 51834

  --1100101001111011    1100101001111100    1100101001111101    1100101001111110    1100101001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51835 - 51839

  --1100101010000000    1100101010000001    1100101010000010    1100101010000011    1100101010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51840 - 51844

  --1100101010000101    1100101010000110    1100101010000111    1100101010001000    1100101010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51845 - 51849

  --1100101010001010    1100101010001011    1100101010001100    1100101010001101    1100101010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51850 - 51854

  --1100101010001111    1100101010010000    1100101010010001    1100101010010010    1100101010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51855 - 51859

  --1100101010010100    1100101010010101    1100101010010110    1100101010010111    1100101010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51860 - 51864

  --1100101010011001    1100101010011010    1100101010011011    1100101010011100    1100101010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51865 - 51869

  --1100101010011110    1100101010011111    1100101010100000    1100101010100001    1100101010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51870 - 51874

  --1100101010100011    1100101010100100    1100101010100101    1100101010100110    1100101010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51875 - 51879

  --1100101010101000    1100101010101001    1100101010101010    1100101010101011    1100101010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51880 - 51884

  --1100101010101101    1100101010101110    1100101010101111    1100101010110000    1100101010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51885 - 51889

  --1100101010110010    1100101010110011    1100101010110100    1100101010110101    1100101010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51890 - 51894

  --1100101010110111    1100101010111000    1100101010111001    1100101010111010    1100101010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51895 - 51899

  --1100101010111100    1100101010111101    1100101010111110    1100101010111111    1100101011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51900 - 51904

  --1100101011000001    1100101011000010    1100101011000011    1100101011000100    1100101011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51905 - 51909

  --1100101011000110    1100101011000111    1100101011001000    1100101011001001    1100101011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51910 - 51914

  --1100101011001011    1100101011001100    1100101011001101    1100101011001110    1100101011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51915 - 51919

  --1100101011010000    1100101011010001    1100101011010010    1100101011010011    1100101011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51920 - 51924

  --1100101011010101    1100101011010110    1100101011010111    1100101011011000    1100101011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51925 - 51929

  --1100101011011010    1100101011011011    1100101011011100    1100101011011101    1100101011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51930 - 51934

  --1100101011011111    1100101011100000    1100101011100001    1100101011100010    1100101011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51935 - 51939

  --1100101011100100    1100101011100101    1100101011100110    1100101011100111    1100101011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51940 - 51944

  --1100101011101001    1100101011101010    1100101011101011    1100101011101100    1100101011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51945 - 51949

  --1100101011101110    1100101011101111    1100101011110000    1100101011110001    1100101011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51950 - 51954

  --1100101011110011    1100101011110100    1100101011110101    1100101011110110    1100101011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51955 - 51959

  --1100101011111000    1100101011111001    1100101011111010    1100101011111011    1100101011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51960 - 51964

  --1100101011111101    1100101011111110    1100101011111111    1100101100000000    1100101100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51965 - 51969

  --1100101100000010    1100101100000011    1100101100000100    1100101100000101    1100101100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51970 - 51974

  --1100101100000111    1100101100001000    1100101100001001    1100101100001010    1100101100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51975 - 51979

  --1100101100001100    1100101100001101    1100101100001110    1100101100001111    1100101100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51980 - 51984

  --1100101100010001    1100101100010010    1100101100010011    1100101100010100    1100101100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51985 - 51989

  --1100101100010110    1100101100010111    1100101100011000    1100101100011001    1100101100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51990 - 51994

  --1100101100011011    1100101100011100    1100101100011101    1100101100011110    1100101100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 51995 - 51999

  --1100101100100000    1100101100100001    1100101100100010    1100101100100011    1100101100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52000 - 52004

  --1100101100100101    1100101100100110    1100101100100111    1100101100101000    1100101100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52005 - 52009

  --1100101100101010    1100101100101011    1100101100101100    1100101100101101    1100101100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52010 - 52014

  --1100101100101111    1100101100110000    1100101100110001    1100101100110010    1100101100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52015 - 52019

  --1100101100110100    1100101100110101    1100101100110110    1100101100110111    1100101100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52020 - 52024

  --1100101100111001    1100101100111010    1100101100111011    1100101100111100    1100101100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52025 - 52029

  --1100101100111110    1100101100111111    1100101101000000    1100101101000001    1100101101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52030 - 52034

  --1100101101000011    1100101101000100    1100101101000101    1100101101000110    1100101101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52035 - 52039

  --1100101101001000    1100101101001001    1100101101001010    1100101101001011    1100101101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52040 - 52044

  --1100101101001101    1100101101001110    1100101101001111    1100101101010000    1100101101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52045 - 52049

  --1100101101010010    1100101101010011    1100101101010100    1100101101010101    1100101101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52050 - 52054

  --1100101101010111    1100101101011000    1100101101011001    1100101101011010    1100101101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52055 - 52059

  --1100101101011100    1100101101011101    1100101101011110    1100101101011111    1100101101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52060 - 52064

  --1100101101100001    1100101101100010    1100101101100011    1100101101100100    1100101101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52065 - 52069

  --1100101101100110    1100101101100111    1100101101101000    1100101101101001    1100101101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52070 - 52074

  --1100101101101011    1100101101101100    1100101101101101    1100101101101110    1100101101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52075 - 52079

  --1100101101110000    1100101101110001    1100101101110010    1100101101110011    1100101101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52080 - 52084

  --1100101101110101    1100101101110110    1100101101110111    1100101101111000    1100101101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52085 - 52089

  --1100101101111010    1100101101111011    1100101101111100    1100101101111101    1100101101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52090 - 52094

  --1100101101111111    1100101110000000    1100101110000001    1100101110000010    1100101110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52095 - 52099

  --1100101110000100    1100101110000101    1100101110000110    1100101110000111    1100101110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52100 - 52104

  --1100101110001001    1100101110001010    1100101110001011    1100101110001100    1100101110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52105 - 52109

  --1100101110001110    1100101110001111    1100101110010000    1100101110010001    1100101110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52110 - 52114

  --1100101110010011    1100101110010100    1100101110010101    1100101110010110    1100101110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52115 - 52119

  --1100101110011000    1100101110011001    1100101110011010    1100101110011011    1100101110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52120 - 52124

  --1100101110011101    1100101110011110    1100101110011111    1100101110100000    1100101110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52125 - 52129

  --1100101110100010    1100101110100011    1100101110100100    1100101110100101    1100101110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52130 - 52134

  --1100101110100111    1100101110101000    1100101110101001    1100101110101010    1100101110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52135 - 52139

  --1100101110101100    1100101110101101    1100101110101110    1100101110101111    1100101110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52140 - 52144

  --1100101110110001    1100101110110010    1100101110110011    1100101110110100    1100101110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52145 - 52149

  --1100101110110110    1100101110110111    1100101110111000    1100101110111001    1100101110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52150 - 52154

  --1100101110111011    1100101110111100    1100101110111101    1100101110111110    1100101110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52155 - 52159

  --1100101111000000    1100101111000001    1100101111000010    1100101111000011    1100101111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52160 - 52164

  --1100101111000101    1100101111000110    1100101111000111    1100101111001000    1100101111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52165 - 52169

  --1100101111001010    1100101111001011    1100101111001100    1100101111001101    1100101111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52170 - 52174

  --1100101111001111    1100101111010000    1100101111010001    1100101111010010    1100101111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52175 - 52179

  --1100101111010100    1100101111010101    1100101111010110    1100101111010111    1100101111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52180 - 52184

  --1100101111011001    1100101111011010    1100101111011011    1100101111011100    1100101111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52185 - 52189

  --1100101111011110    1100101111011111    1100101111100000    1100101111100001    1100101111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52190 - 52194

  --1100101111100011    1100101111100100    1100101111100101    1100101111100110    1100101111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52195 - 52199

  --1100101111101000    1100101111101001    1100101111101010    1100101111101011    1100101111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52200 - 52204

  --1100101111101101    1100101111101110    1100101111101111    1100101111110000    1100101111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52205 - 52209

  --1100101111110010    1100101111110011    1100101111110100    1100101111110101    1100101111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52210 - 52214

  --1100101111110111    1100101111111000    1100101111111001    1100101111111010    1100101111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52215 - 52219

  --1100101111111100    1100101111111101    1100101111111110    1100101111111111    1100110000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52220 - 52224

  --1100110000000001    1100110000000010    1100110000000011    1100110000000100    1100110000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52225 - 52229

  --1100110000000110    1100110000000111    1100110000001000    1100110000001001    1100110000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52230 - 52234

  --1100110000001011    1100110000001100    1100110000001101    1100110000001110    1100110000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52235 - 52239

  --1100110000010000    1100110000010001    1100110000010010    1100110000010011    1100110000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52240 - 52244

  --1100110000010101    1100110000010110    1100110000010111    1100110000011000    1100110000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52245 - 52249

  --1100110000011010    1100110000011011    1100110000011100    1100110000011101    1100110000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52250 - 52254

  --1100110000011111    1100110000100000    1100110000100001    1100110000100010    1100110000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52255 - 52259

  --1100110000100100    1100110000100101    1100110000100110    1100110000100111    1100110000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52260 - 52264

  --1100110000101001    1100110000101010    1100110000101011    1100110000101100    1100110000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52265 - 52269

  --1100110000101110    1100110000101111    1100110000110000    1100110000110001    1100110000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52270 - 52274

  --1100110000110011    1100110000110100    1100110000110101    1100110000110110    1100110000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52275 - 52279

  --1100110000111000    1100110000111001    1100110000111010    1100110000111011    1100110000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52280 - 52284

  --1100110000111101    1100110000111110    1100110000111111    1100110001000000    1100110001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52285 - 52289

  --1100110001000010    1100110001000011    1100110001000100    1100110001000101    1100110001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52290 - 52294

  --1100110001000111    1100110001001000    1100110001001001    1100110001001010    1100110001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52295 - 52299

  --1100110001001100    1100110001001101    1100110001001110    1100110001001111    1100110001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52300 - 52304

  --1100110001010001    1100110001010010    1100110001010011    1100110001010100    1100110001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52305 - 52309

  --1100110001010110    1100110001010111    1100110001011000    1100110001011001    1100110001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52310 - 52314

  --1100110001011011    1100110001011100    1100110001011101    1100110001011110    1100110001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52315 - 52319

  --1100110001100000    1100110001100001    1100110001100010    1100110001100011    1100110001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52320 - 52324

  --1100110001100101    1100110001100110    1100110001100111    1100110001101000    1100110001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52325 - 52329

  --1100110001101010    1100110001101011    1100110001101100    1100110001101101    1100110001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52330 - 52334

  --1100110001101111    1100110001110000    1100110001110001    1100110001110010    1100110001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52335 - 52339

  --1100110001110100    1100110001110101    1100110001110110    1100110001110111    1100110001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52340 - 52344

  --1100110001111001    1100110001111010    1100110001111011    1100110001111100    1100110001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52345 - 52349

  --1100110001111110    1100110001111111    1100110010000000    1100110010000001    1100110010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52350 - 52354

  --1100110010000011    1100110010000100    1100110010000101    1100110010000110    1100110010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52355 - 52359

  --1100110010001000    1100110010001001    1100110010001010    1100110010001011    1100110010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52360 - 52364

  --1100110010001101    1100110010001110    1100110010001111    1100110010010000    1100110010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52365 - 52369

  --1100110010010010    1100110010010011    1100110010010100    1100110010010101    1100110010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52370 - 52374

  --1100110010010111    1100110010011000    1100110010011001    1100110010011010    1100110010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52375 - 52379

  --1100110010011100    1100110010011101    1100110010011110    1100110010011111    1100110010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52380 - 52384

  --1100110010100001    1100110010100010    1100110010100011    1100110010100100    1100110010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52385 - 52389

  --1100110010100110    1100110010100111    1100110010101000    1100110010101001    1100110010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52390 - 52394

  --1100110010101011    1100110010101100    1100110010101101    1100110010101110    1100110010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52395 - 52399

  --1100110010110000    1100110010110001    1100110010110010    1100110010110011    1100110010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52400 - 52404

  --1100110010110101    1100110010110110    1100110010110111    1100110010111000    1100110010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52405 - 52409

  --1100110010111010    1100110010111011    1100110010111100    1100110010111101    1100110010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52410 - 52414

  --1100110010111111    1100110011000000    1100110011000001    1100110011000010    1100110011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52415 - 52419

  --1100110011000100    1100110011000101    1100110011000110    1100110011000111    1100110011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52420 - 52424

  --1100110011001001    1100110011001010    1100110011001011    1100110011001100    1100110011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52425 - 52429

  --1100110011001110    1100110011001111    1100110011010000    1100110011010001    1100110011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52430 - 52434

  --1100110011010011    1100110011010100    1100110011010101    1100110011010110    1100110011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52435 - 52439

  --1100110011011000    1100110011011001    1100110011011010    1100110011011011    1100110011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52440 - 52444

  --1100110011011101    1100110011011110    1100110011011111    1100110011100000    1100110011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52445 - 52449

  --1100110011100010    1100110011100011    1100110011100100    1100110011100101    1100110011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52450 - 52454

  --1100110011100111    1100110011101000    1100110011101001    1100110011101010    1100110011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52455 - 52459

  --1100110011101100    1100110011101101    1100110011101110    1100110011101111    1100110011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52460 - 52464

  --1100110011110001    1100110011110010    1100110011110011    1100110011110100    1100110011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52465 - 52469

  --1100110011110110    1100110011110111    1100110011111000    1100110011111001    1100110011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52470 - 52474

  --1100110011111011    1100110011111100    1100110011111101    1100110011111110    1100110011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52475 - 52479

  --1100110100000000    1100110100000001    1100110100000010    1100110100000011    1100110100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52480 - 52484

  --1100110100000101    1100110100000110    1100110100000111    1100110100001000    1100110100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52485 - 52489

  --1100110100001010    1100110100001011    1100110100001100    1100110100001101    1100110100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52490 - 52494

  --1100110100001111    1100110100010000    1100110100010001    1100110100010010    1100110100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52495 - 52499

  --1100110100010100    1100110100010101    1100110100010110    1100110100010111    1100110100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52500 - 52504

  --1100110100011001    1100110100011010    1100110100011011    1100110100011100    1100110100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52505 - 52509

  --1100110100011110    1100110100011111    1100110100100000    1100110100100001    1100110100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52510 - 52514

  --1100110100100011    1100110100100100    1100110100100101    1100110100100110    1100110100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52515 - 52519

  --1100110100101000    1100110100101001    1100110100101010    1100110100101011    1100110100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52520 - 52524

  --1100110100101101    1100110100101110    1100110100101111    1100110100110000    1100110100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52525 - 52529

  --1100110100110010    1100110100110011    1100110100110100    1100110100110101    1100110100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52530 - 52534

  --1100110100110111    1100110100111000    1100110100111001    1100110100111010    1100110100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52535 - 52539

  --1100110100111100    1100110100111101    1100110100111110    1100110100111111    1100110101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52540 - 52544

  --1100110101000001    1100110101000010    1100110101000011    1100110101000100    1100110101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52545 - 52549

  --1100110101000110    1100110101000111    1100110101001000    1100110101001001    1100110101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52550 - 52554

  --1100110101001011    1100110101001100    1100110101001101    1100110101001110    1100110101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52555 - 52559

  --1100110101010000    1100110101010001    1100110101010010    1100110101010011    1100110101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52560 - 52564

  --1100110101010101    1100110101010110    1100110101010111    1100110101011000    1100110101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52565 - 52569

  --1100110101011010    1100110101011011    1100110101011100    1100110101011101    1100110101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52570 - 52574

  --1100110101011111    1100110101100000    1100110101100001    1100110101100010    1100110101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52575 - 52579

  --1100110101100100    1100110101100101    1100110101100110    1100110101100111    1100110101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52580 - 52584

  --1100110101101001    1100110101101010    1100110101101011    1100110101101100    1100110101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52585 - 52589

  --1100110101101110    1100110101101111    1100110101110000    1100110101110001    1100110101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52590 - 52594

  --1100110101110011    1100110101110100    1100110101110101    1100110101110110    1100110101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52595 - 52599

  --1100110101111000    1100110101111001    1100110101111010    1100110101111011    1100110101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52600 - 52604

  --1100110101111101    1100110101111110    1100110101111111    1100110110000000    1100110110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52605 - 52609

  --1100110110000010    1100110110000011    1100110110000100    1100110110000101    1100110110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52610 - 52614

  --1100110110000111    1100110110001000    1100110110001001    1100110110001010    1100110110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52615 - 52619

  --1100110110001100    1100110110001101    1100110110001110    1100110110001111    1100110110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52620 - 52624

  --1100110110010001    1100110110010010    1100110110010011    1100110110010100    1100110110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52625 - 52629

  --1100110110010110    1100110110010111    1100110110011000    1100110110011001    1100110110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52630 - 52634

  --1100110110011011    1100110110011100    1100110110011101    1100110110011110    1100110110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52635 - 52639

  --1100110110100000    1100110110100001    1100110110100010    1100110110100011    1100110110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52640 - 52644

  --1100110110100101    1100110110100110    1100110110100111    1100110110101000    1100110110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52645 - 52649

  --1100110110101010    1100110110101011    1100110110101100    1100110110101101    1100110110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52650 - 52654

  --1100110110101111    1100110110110000    1100110110110001    1100110110110010    1100110110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52655 - 52659

  --1100110110110100    1100110110110101    1100110110110110    1100110110110111    1100110110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52660 - 52664

  --1100110110111001    1100110110111010    1100110110111011    1100110110111100    1100110110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52665 - 52669

  --1100110110111110    1100110110111111    1100110111000000    1100110111000001    1100110111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52670 - 52674

  --1100110111000011    1100110111000100    1100110111000101    1100110111000110    1100110111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52675 - 52679

  --1100110111001000    1100110111001001    1100110111001010    1100110111001011    1100110111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52680 - 52684

  --1100110111001101    1100110111001110    1100110111001111    1100110111010000    1100110111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52685 - 52689

  --1100110111010010    1100110111010011    1100110111010100    1100110111010101    1100110111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52690 - 52694

  --1100110111010111    1100110111011000    1100110111011001    1100110111011010    1100110111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52695 - 52699

  --1100110111011100    1100110111011101    1100110111011110    1100110111011111    1100110111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52700 - 52704

  --1100110111100001    1100110111100010    1100110111100011    1100110111100100    1100110111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52705 - 52709

  --1100110111100110    1100110111100111    1100110111101000    1100110111101001    1100110111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52710 - 52714

  --1100110111101011    1100110111101100    1100110111101101    1100110111101110    1100110111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52715 - 52719

  --1100110111110000    1100110111110001    1100110111110010    1100110111110011    1100110111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52720 - 52724

  --1100110111110101    1100110111110110    1100110111110111    1100110111111000    1100110111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52725 - 52729

  --1100110111111010    1100110111111011    1100110111111100    1100110111111101    1100110111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52730 - 52734

  --1100110111111111    1100111000000000    1100111000000001    1100111000000010    1100111000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52735 - 52739

  --1100111000000100    1100111000000101    1100111000000110    1100111000000111    1100111000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52740 - 52744

  --1100111000001001    1100111000001010    1100111000001011    1100111000001100    1100111000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52745 - 52749

  --1100111000001110    1100111000001111    1100111000010000    1100111000010001    1100111000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52750 - 52754

  --1100111000010011    1100111000010100    1100111000010101    1100111000010110    1100111000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52755 - 52759

  --1100111000011000    1100111000011001    1100111000011010    1100111000011011    1100111000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52760 - 52764

  --1100111000011101    1100111000011110    1100111000011111    1100111000100000    1100111000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52765 - 52769

  --1100111000100010    1100111000100011    1100111000100100    1100111000100101    1100111000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52770 - 52774

  --1100111000100111    1100111000101000    1100111000101001    1100111000101010    1100111000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52775 - 52779

  --1100111000101100    1100111000101101    1100111000101110    1100111000101111    1100111000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52780 - 52784

  --1100111000110001    1100111000110010    1100111000110011    1100111000110100    1100111000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52785 - 52789

  --1100111000110110    1100111000110111    1100111000111000    1100111000111001    1100111000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52790 - 52794

  --1100111000111011    1100111000111100    1100111000111101    1100111000111110    1100111000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52795 - 52799

  --1100111001000000    1100111001000001    1100111001000010    1100111001000011    1100111001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52800 - 52804

  --1100111001000101    1100111001000110    1100111001000111    1100111001001000    1100111001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52805 - 52809

  --1100111001001010    1100111001001011    1100111001001100    1100111001001101    1100111001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52810 - 52814

  --1100111001001111    1100111001010000    1100111001010001    1100111001010010    1100111001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52815 - 52819

  --1100111001010100    1100111001010101    1100111001010110    1100111001010111    1100111001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52820 - 52824

  --1100111001011001    1100111001011010    1100111001011011    1100111001011100    1100111001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52825 - 52829

  --1100111001011110    1100111001011111    1100111001100000    1100111001100001    1100111001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52830 - 52834

  --1100111001100011    1100111001100100    1100111001100101    1100111001100110    1100111001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52835 - 52839

  --1100111001101000    1100111001101001    1100111001101010    1100111001101011    1100111001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52840 - 52844

  --1100111001101101    1100111001101110    1100111001101111    1100111001110000    1100111001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52845 - 52849

  --1100111001110010    1100111001110011    1100111001110100    1100111001110101    1100111001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52850 - 52854

  --1100111001110111    1100111001111000    1100111001111001    1100111001111010    1100111001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52855 - 52859

  --1100111001111100    1100111001111101    1100111001111110    1100111001111111    1100111010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52860 - 52864

  --1100111010000001    1100111010000010    1100111010000011    1100111010000100    1100111010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52865 - 52869

  --1100111010000110    1100111010000111    1100111010001000    1100111010001001    1100111010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52870 - 52874

  --1100111010001011    1100111010001100    1100111010001101    1100111010001110    1100111010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52875 - 52879

  --1100111010010000    1100111010010001    1100111010010010    1100111010010011    1100111010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52880 - 52884

  --1100111010010101    1100111010010110    1100111010010111    1100111010011000    1100111010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52885 - 52889

  --1100111010011010    1100111010011011    1100111010011100    1100111010011101    1100111010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52890 - 52894

  --1100111010011111    1100111010100000    1100111010100001    1100111010100010    1100111010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52895 - 52899

  --1100111010100100    1100111010100101    1100111010100110    1100111010100111    1100111010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52900 - 52904

  --1100111010101001    1100111010101010    1100111010101011    1100111010101100    1100111010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52905 - 52909

  --1100111010101110    1100111010101111    1100111010110000    1100111010110001    1100111010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52910 - 52914

  --1100111010110011    1100111010110100    1100111010110101    1100111010110110    1100111010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52915 - 52919

  --1100111010111000    1100111010111001    1100111010111010    1100111010111011    1100111010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52920 - 52924

  --1100111010111101    1100111010111110    1100111010111111    1100111011000000    1100111011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52925 - 52929

  --1100111011000010    1100111011000011    1100111011000100    1100111011000101    1100111011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52930 - 52934

  --1100111011000111    1100111011001000    1100111011001001    1100111011001010    1100111011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52935 - 52939

  --1100111011001100    1100111011001101    1100111011001110    1100111011001111    1100111011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52940 - 52944

  --1100111011010001    1100111011010010    1100111011010011    1100111011010100    1100111011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52945 - 52949

  --1100111011010110    1100111011010111    1100111011011000    1100111011011001    1100111011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52950 - 52954

  --1100111011011011    1100111011011100    1100111011011101    1100111011011110    1100111011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52955 - 52959

  --1100111011100000    1100111011100001    1100111011100010    1100111011100011    1100111011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52960 - 52964

  --1100111011100101    1100111011100110    1100111011100111    1100111011101000    1100111011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52965 - 52969

  --1100111011101010    1100111011101011    1100111011101100    1100111011101101    1100111011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52970 - 52974

  --1100111011101111    1100111011110000    1100111011110001    1100111011110010    1100111011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52975 - 52979

  --1100111011110100    1100111011110101    1100111011110110    1100111011110111    1100111011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52980 - 52984

  --1100111011111001    1100111011111010    1100111011111011    1100111011111100    1100111011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52985 - 52989

  --1100111011111110    1100111011111111    1100111100000000    1100111100000001    1100111100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52990 - 52994

  --1100111100000011    1100111100000100    1100111100000101    1100111100000110    1100111100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 52995 - 52999

  --1100111100001000    1100111100001001    1100111100001010    1100111100001011    1100111100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53000 - 53004

  --1100111100001101    1100111100001110    1100111100001111    1100111100010000    1100111100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53005 - 53009

  --1100111100010010    1100111100010011    1100111100010100    1100111100010101    1100111100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53010 - 53014

  --1100111100010111    1100111100011000    1100111100011001    1100111100011010    1100111100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53015 - 53019

  --1100111100011100    1100111100011101    1100111100011110    1100111100011111    1100111100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53020 - 53024

  --1100111100100001    1100111100100010    1100111100100011    1100111100100100    1100111100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53025 - 53029

  --1100111100100110    1100111100100111    1100111100101000    1100111100101001    1100111100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53030 - 53034

  --1100111100101011    1100111100101100    1100111100101101    1100111100101110    1100111100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53035 - 53039

  --1100111100110000    1100111100110001    1100111100110010    1100111100110011    1100111100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53040 - 53044

  --1100111100110101    1100111100110110    1100111100110111    1100111100111000    1100111100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53045 - 53049

  --1100111100111010    1100111100111011    1100111100111100    1100111100111101    1100111100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53050 - 53054

  --1100111100111111    1100111101000000    1100111101000001    1100111101000010    1100111101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53055 - 53059

  --1100111101000100    1100111101000101    1100111101000110    1100111101000111    1100111101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53060 - 53064

  --1100111101001001    1100111101001010    1100111101001011    1100111101001100    1100111101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53065 - 53069

  --1100111101001110    1100111101001111    1100111101010000    1100111101010001    1100111101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53070 - 53074

  --1100111101010011    1100111101010100    1100111101010101    1100111101010110    1100111101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53075 - 53079

  --1100111101011000    1100111101011001    1100111101011010    1100111101011011    1100111101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53080 - 53084

  --1100111101011101    1100111101011110    1100111101011111    1100111101100000    1100111101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53085 - 53089

  --1100111101100010    1100111101100011    1100111101100100    1100111101100101    1100111101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53090 - 53094

  --1100111101100111    1100111101101000    1100111101101001    1100111101101010    1100111101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53095 - 53099

  --1100111101101100    1100111101101101    1100111101101110    1100111101101111    1100111101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53100 - 53104

  --1100111101110001    1100111101110010    1100111101110011    1100111101110100    1100111101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53105 - 53109

  --1100111101110110    1100111101110111    1100111101111000    1100111101111001    1100111101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53110 - 53114

  --1100111101111011    1100111101111100    1100111101111101    1100111101111110    1100111101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53115 - 53119

  --1100111110000000    1100111110000001    1100111110000010    1100111110000011    1100111110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53120 - 53124

  --1100111110000101    1100111110000110    1100111110000111    1100111110001000    1100111110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53125 - 53129

  --1100111110001010    1100111110001011    1100111110001100    1100111110001101    1100111110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53130 - 53134

  --1100111110001111    1100111110010000    1100111110010001    1100111110010010    1100111110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53135 - 53139

  --1100111110010100    1100111110010101    1100111110010110    1100111110010111    1100111110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53140 - 53144

  --1100111110011001    1100111110011010    1100111110011011    1100111110011100    1100111110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53145 - 53149

  --1100111110011110    1100111110011111    1100111110100000    1100111110100001    1100111110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53150 - 53154

  --1100111110100011    1100111110100100    1100111110100101    1100111110100110    1100111110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53155 - 53159

  --1100111110101000    1100111110101001    1100111110101010    1100111110101011    1100111110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53160 - 53164

  --1100111110101101    1100111110101110    1100111110101111    1100111110110000    1100111110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53165 - 53169

  --1100111110110010    1100111110110011    1100111110110100    1100111110110101    1100111110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53170 - 53174

  --1100111110110111    1100111110111000    1100111110111001    1100111110111010    1100111110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53175 - 53179

  --1100111110111100    1100111110111101    1100111110111110    1100111110111111    1100111111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53180 - 53184

  --1100111111000001    1100111111000010    1100111111000011    1100111111000100    1100111111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53185 - 53189

  --1100111111000110    1100111111000111    1100111111001000    1100111111001001    1100111111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53190 - 53194

  --1100111111001011    1100111111001100    1100111111001101    1100111111001110    1100111111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53195 - 53199

  --1100111111010000    1100111111010001    1100111111010010    1100111111010011    1100111111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53200 - 53204

  --1100111111010101    1100111111010110    1100111111010111    1100111111011000    1100111111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53205 - 53209

  --1100111111011010    1100111111011011    1100111111011100    1100111111011101    1100111111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53210 - 53214

  --1100111111011111    1100111111100000    1100111111100001    1100111111100010    1100111111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53215 - 53219

  --1100111111100100    1100111111100101    1100111111100110    1100111111100111    1100111111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53220 - 53224

  --1100111111101001    1100111111101010    1100111111101011    1100111111101100    1100111111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53225 - 53229

  --1100111111101110    1100111111101111    1100111111110000    1100111111110001    1100111111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53230 - 53234

  --1100111111110011    1100111111110100    1100111111110101    1100111111110110    1100111111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53235 - 53239

  --1100111111111000    1100111111111001    1100111111111010    1100111111111011    1100111111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53240 - 53244

  --1100111111111101    1100111111111110    1100111111111111    1101000000000000    1101000000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53245 - 53249

  --1101000000000010    1101000000000011    1101000000000100    1101000000000101    1101000000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53250 - 53254

  --1101000000000111    1101000000001000    1101000000001001    1101000000001010    1101000000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53255 - 53259

  --1101000000001100    1101000000001101    1101000000001110    1101000000001111    1101000000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53260 - 53264

  --1101000000010001    1101000000010010    1101000000010011    1101000000010100    1101000000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53265 - 53269

  --1101000000010110    1101000000010111    1101000000011000    1101000000011001    1101000000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53270 - 53274

  --1101000000011011    1101000000011100    1101000000011101    1101000000011110    1101000000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53275 - 53279

  --1101000000100000    1101000000100001    1101000000100010    1101000000100011    1101000000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53280 - 53284

  --1101000000100101    1101000000100110    1101000000100111    1101000000101000    1101000000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53285 - 53289

  --1101000000101010    1101000000101011    1101000000101100    1101000000101101    1101000000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53290 - 53294

  --1101000000101111    1101000000110000    1101000000110001    1101000000110010    1101000000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53295 - 53299

  --1101000000110100    1101000000110101    1101000000110110    1101000000110111    1101000000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53300 - 53304

  --1101000000111001    1101000000111010    1101000000111011    1101000000111100    1101000000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53305 - 53309

  --1101000000111110    1101000000111111    1101000001000000    1101000001000001    1101000001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53310 - 53314

  --1101000001000011    1101000001000100    1101000001000101    1101000001000110    1101000001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53315 - 53319

  --1101000001001000    1101000001001001    1101000001001010    1101000001001011    1101000001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53320 - 53324

  --1101000001001101    1101000001001110    1101000001001111    1101000001010000    1101000001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53325 - 53329

  --1101000001010010    1101000001010011    1101000001010100    1101000001010101    1101000001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53330 - 53334

  --1101000001010111    1101000001011000    1101000001011001    1101000001011010    1101000001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53335 - 53339

  --1101000001011100    1101000001011101    1101000001011110    1101000001011111    1101000001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53340 - 53344

  --1101000001100001    1101000001100010    1101000001100011    1101000001100100    1101000001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53345 - 53349

  --1101000001100110    1101000001100111    1101000001101000    1101000001101001    1101000001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53350 - 53354

  --1101000001101011    1101000001101100    1101000001101101    1101000001101110    1101000001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53355 - 53359

  --1101000001110000    1101000001110001    1101000001110010    1101000001110011    1101000001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53360 - 53364

  --1101000001110101    1101000001110110    1101000001110111    1101000001111000    1101000001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53365 - 53369

  --1101000001111010    1101000001111011    1101000001111100    1101000001111101    1101000001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53370 - 53374

  --1101000001111111    1101000010000000    1101000010000001    1101000010000010    1101000010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53375 - 53379

  --1101000010000100    1101000010000101    1101000010000110    1101000010000111    1101000010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53380 - 53384

  --1101000010001001    1101000010001010    1101000010001011    1101000010001100    1101000010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53385 - 53389

  --1101000010001110    1101000010001111    1101000010010000    1101000010010001    1101000010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53390 - 53394

  --1101000010010011    1101000010010100    1101000010010101    1101000010010110    1101000010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53395 - 53399

  --1101000010011000    1101000010011001    1101000010011010    1101000010011011    1101000010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53400 - 53404

  --1101000010011101    1101000010011110    1101000010011111    1101000010100000    1101000010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53405 - 53409

  --1101000010100010    1101000010100011    1101000010100100    1101000010100101    1101000010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53410 - 53414

  --1101000010100111    1101000010101000    1101000010101001    1101000010101010    1101000010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53415 - 53419

  --1101000010101100    1101000010101101    1101000010101110    1101000010101111    1101000010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53420 - 53424

  --1101000010110001    1101000010110010    1101000010110011    1101000010110100    1101000010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53425 - 53429

  --1101000010110110    1101000010110111    1101000010111000    1101000010111001    1101000010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53430 - 53434

  --1101000010111011    1101000010111100    1101000010111101    1101000010111110    1101000010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53435 - 53439

  --1101000011000000    1101000011000001    1101000011000010    1101000011000011    1101000011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53440 - 53444

  --1101000011000101    1101000011000110    1101000011000111    1101000011001000    1101000011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53445 - 53449

  --1101000011001010    1101000011001011    1101000011001100    1101000011001101    1101000011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53450 - 53454

  --1101000011001111    1101000011010000    1101000011010001    1101000011010010    1101000011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53455 - 53459

  --1101000011010100    1101000011010101    1101000011010110    1101000011010111    1101000011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53460 - 53464

  --1101000011011001    1101000011011010    1101000011011011    1101000011011100    1101000011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53465 - 53469

  --1101000011011110    1101000011011111    1101000011100000    1101000011100001    1101000011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53470 - 53474

  --1101000011100011    1101000011100100    1101000011100101    1101000011100110    1101000011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53475 - 53479

  --1101000011101000    1101000011101001    1101000011101010    1101000011101011    1101000011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53480 - 53484

  --1101000011101101    1101000011101110    1101000011101111    1101000011110000    1101000011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53485 - 53489

  --1101000011110010    1101000011110011    1101000011110100    1101000011110101    1101000011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53490 - 53494

  --1101000011110111    1101000011111000    1101000011111001    1101000011111010    1101000011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53495 - 53499

  --1101000011111100    1101000011111101    1101000011111110    1101000011111111    1101000100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53500 - 53504

  --1101000100000001    1101000100000010    1101000100000011    1101000100000100    1101000100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53505 - 53509

  --1101000100000110    1101000100000111    1101000100001000    1101000100001001    1101000100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53510 - 53514

  --1101000100001011    1101000100001100    1101000100001101    1101000100001110    1101000100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53515 - 53519

  --1101000100010000    1101000100010001    1101000100010010    1101000100010011    1101000100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53520 - 53524

  --1101000100010101    1101000100010110    1101000100010111    1101000100011000    1101000100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53525 - 53529

  --1101000100011010    1101000100011011    1101000100011100    1101000100011101    1101000100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53530 - 53534

  --1101000100011111    1101000100100000    1101000100100001    1101000100100010    1101000100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53535 - 53539

  --1101000100100100    1101000100100101    1101000100100110    1101000100100111    1101000100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53540 - 53544

  --1101000100101001    1101000100101010    1101000100101011    1101000100101100    1101000100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53545 - 53549

  --1101000100101110    1101000100101111    1101000100110000    1101000100110001    1101000100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53550 - 53554

  --1101000100110011    1101000100110100    1101000100110101    1101000100110110    1101000100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53555 - 53559

  --1101000100111000    1101000100111001    1101000100111010    1101000100111011    1101000100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53560 - 53564

  --1101000100111101    1101000100111110    1101000100111111    1101000101000000    1101000101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53565 - 53569

  --1101000101000010    1101000101000011    1101000101000100    1101000101000101    1101000101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53570 - 53574

  --1101000101000111    1101000101001000    1101000101001001    1101000101001010    1101000101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53575 - 53579

  --1101000101001100    1101000101001101    1101000101001110    1101000101001111    1101000101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53580 - 53584

  --1101000101010001    1101000101010010    1101000101010011    1101000101010100    1101000101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53585 - 53589

  --1101000101010110    1101000101010111    1101000101011000    1101000101011001    1101000101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53590 - 53594

  --1101000101011011    1101000101011100    1101000101011101    1101000101011110    1101000101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53595 - 53599

  --1101000101100000    1101000101100001    1101000101100010    1101000101100011    1101000101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53600 - 53604

  --1101000101100101    1101000101100110    1101000101100111    1101000101101000    1101000101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53605 - 53609

  --1101000101101010    1101000101101011    1101000101101100    1101000101101101    1101000101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53610 - 53614

  --1101000101101111    1101000101110000    1101000101110001    1101000101110010    1101000101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53615 - 53619

  --1101000101110100    1101000101110101    1101000101110110    1101000101110111    1101000101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53620 - 53624

  --1101000101111001    1101000101111010    1101000101111011    1101000101111100    1101000101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53625 - 53629

  --1101000101111110    1101000101111111    1101000110000000    1101000110000001    1101000110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53630 - 53634

  --1101000110000011    1101000110000100    1101000110000101    1101000110000110    1101000110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53635 - 53639

  --1101000110001000    1101000110001001    1101000110001010    1101000110001011    1101000110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53640 - 53644

  --1101000110001101    1101000110001110    1101000110001111    1101000110010000    1101000110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53645 - 53649

  --1101000110010010    1101000110010011    1101000110010100    1101000110010101    1101000110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53650 - 53654

  --1101000110010111    1101000110011000    1101000110011001    1101000110011010    1101000110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53655 - 53659

  --1101000110011100    1101000110011101    1101000110011110    1101000110011111    1101000110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53660 - 53664

  --1101000110100001    1101000110100010    1101000110100011    1101000110100100    1101000110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53665 - 53669

  --1101000110100110    1101000110100111    1101000110101000    1101000110101001    1101000110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53670 - 53674

  --1101000110101011    1101000110101100    1101000110101101    1101000110101110    1101000110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53675 - 53679

  --1101000110110000    1101000110110001    1101000110110010    1101000110110011    1101000110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53680 - 53684

  --1101000110110101    1101000110110110    1101000110110111    1101000110111000    1101000110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53685 - 53689

  --1101000110111010    1101000110111011    1101000110111100    1101000110111101    1101000110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53690 - 53694

  --1101000110111111    1101000111000000    1101000111000001    1101000111000010    1101000111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53695 - 53699

  --1101000111000100    1101000111000101    1101000111000110    1101000111000111    1101000111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53700 - 53704

  --1101000111001001    1101000111001010    1101000111001011    1101000111001100    1101000111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53705 - 53709

  --1101000111001110    1101000111001111    1101000111010000    1101000111010001    1101000111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53710 - 53714

  --1101000111010011    1101000111010100    1101000111010101    1101000111010110    1101000111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53715 - 53719

  --1101000111011000    1101000111011001    1101000111011010    1101000111011011    1101000111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53720 - 53724

  --1101000111011101    1101000111011110    1101000111011111    1101000111100000    1101000111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53725 - 53729

  --1101000111100010    1101000111100011    1101000111100100    1101000111100101    1101000111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53730 - 53734

  --1101000111100111    1101000111101000    1101000111101001    1101000111101010    1101000111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53735 - 53739

  --1101000111101100    1101000111101101    1101000111101110    1101000111101111    1101000111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53740 - 53744

  --1101000111110001    1101000111110010    1101000111110011    1101000111110100    1101000111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53745 - 53749

  --1101000111110110    1101000111110111    1101000111111000    1101000111111001    1101000111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53750 - 53754

  --1101000111111011    1101000111111100    1101000111111101    1101000111111110    1101000111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53755 - 53759

  --1101001000000000    1101001000000001    1101001000000010    1101001000000011    1101001000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53760 - 53764

  --1101001000000101    1101001000000110    1101001000000111    1101001000001000    1101001000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53765 - 53769

  --1101001000001010    1101001000001011    1101001000001100    1101001000001101    1101001000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53770 - 53774

  --1101001000001111    1101001000010000    1101001000010001    1101001000010010    1101001000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53775 - 53779

  --1101001000010100    1101001000010101    1101001000010110    1101001000010111    1101001000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53780 - 53784

  --1101001000011001    1101001000011010    1101001000011011    1101001000011100    1101001000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53785 - 53789

  --1101001000011110    1101001000011111    1101001000100000    1101001000100001    1101001000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53790 - 53794

  --1101001000100011    1101001000100100    1101001000100101    1101001000100110    1101001000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53795 - 53799

  --1101001000101000    1101001000101001    1101001000101010    1101001000101011    1101001000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53800 - 53804

  --1101001000101101    1101001000101110    1101001000101111    1101001000110000    1101001000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53805 - 53809

  --1101001000110010    1101001000110011    1101001000110100    1101001000110101    1101001000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53810 - 53814

  --1101001000110111    1101001000111000    1101001000111001    1101001000111010    1101001000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53815 - 53819

  --1101001000111100    1101001000111101    1101001000111110    1101001000111111    1101001001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53820 - 53824

  --1101001001000001    1101001001000010    1101001001000011    1101001001000100    1101001001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53825 - 53829

  --1101001001000110    1101001001000111    1101001001001000    1101001001001001    1101001001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53830 - 53834

  --1101001001001011    1101001001001100    1101001001001101    1101001001001110    1101001001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53835 - 53839

  --1101001001010000    1101001001010001    1101001001010010    1101001001010011    1101001001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53840 - 53844

  --1101001001010101    1101001001010110    1101001001010111    1101001001011000    1101001001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53845 - 53849

  --1101001001011010    1101001001011011    1101001001011100    1101001001011101    1101001001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53850 - 53854

  --1101001001011111    1101001001100000    1101001001100001    1101001001100010    1101001001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53855 - 53859

  --1101001001100100    1101001001100101    1101001001100110    1101001001100111    1101001001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53860 - 53864

  --1101001001101001    1101001001101010    1101001001101011    1101001001101100    1101001001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53865 - 53869

  --1101001001101110    1101001001101111    1101001001110000    1101001001110001    1101001001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53870 - 53874

  --1101001001110011    1101001001110100    1101001001110101    1101001001110110    1101001001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53875 - 53879

  --1101001001111000    1101001001111001    1101001001111010    1101001001111011    1101001001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53880 - 53884

  --1101001001111101    1101001001111110    1101001001111111    1101001010000000    1101001010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53885 - 53889

  --1101001010000010    1101001010000011    1101001010000100    1101001010000101    1101001010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53890 - 53894

  --1101001010000111    1101001010001000    1101001010001001    1101001010001010    1101001010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53895 - 53899

  --1101001010001100    1101001010001101    1101001010001110    1101001010001111    1101001010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53900 - 53904

  --1101001010010001    1101001010010010    1101001010010011    1101001010010100    1101001010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53905 - 53909

  --1101001010010110    1101001010010111    1101001010011000    1101001010011001    1101001010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53910 - 53914

  --1101001010011011    1101001010011100    1101001010011101    1101001010011110    1101001010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53915 - 53919

  --1101001010100000    1101001010100001    1101001010100010    1101001010100011    1101001010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53920 - 53924

  --1101001010100101    1101001010100110    1101001010100111    1101001010101000    1101001010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53925 - 53929

  --1101001010101010    1101001010101011    1101001010101100    1101001010101101    1101001010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53930 - 53934

  --1101001010101111    1101001010110000    1101001010110001    1101001010110010    1101001010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53935 - 53939

  --1101001010110100    1101001010110101    1101001010110110    1101001010110111    1101001010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53940 - 53944

  --1101001010111001    1101001010111010    1101001010111011    1101001010111100    1101001010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53945 - 53949

  --1101001010111110    1101001010111111    1101001011000000    1101001011000001    1101001011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53950 - 53954

  --1101001011000011    1101001011000100    1101001011000101    1101001011000110    1101001011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53955 - 53959

  --1101001011001000    1101001011001001    1101001011001010    1101001011001011    1101001011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53960 - 53964

  --1101001011001101    1101001011001110    1101001011001111    1101001011010000    1101001011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53965 - 53969

  --1101001011010010    1101001011010011    1101001011010100    1101001011010101    1101001011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53970 - 53974

  --1101001011010111    1101001011011000    1101001011011001    1101001011011010    1101001011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53975 - 53979

  --1101001011011100    1101001011011101    1101001011011110    1101001011011111    1101001011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53980 - 53984

  --1101001011100001    1101001011100010    1101001011100011    1101001011100100    1101001011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53985 - 53989

  --1101001011100110    1101001011100111    1101001011101000    1101001011101001    1101001011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53990 - 53994

  --1101001011101011    1101001011101100    1101001011101101    1101001011101110    1101001011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 53995 - 53999

  --1101001011110000    1101001011110001    1101001011110010    1101001011110011    1101001011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54000 - 54004

  --1101001011110101    1101001011110110    1101001011110111    1101001011111000    1101001011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54005 - 54009

  --1101001011111010    1101001011111011    1101001011111100    1101001011111101    1101001011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54010 - 54014

  --1101001011111111    1101001100000000    1101001100000001    1101001100000010    1101001100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54015 - 54019

  --1101001100000100    1101001100000101    1101001100000110    1101001100000111    1101001100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54020 - 54024

  --1101001100001001    1101001100001010    1101001100001011    1101001100001100    1101001100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54025 - 54029

  --1101001100001110    1101001100001111    1101001100010000    1101001100010001    1101001100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54030 - 54034

  --1101001100010011    1101001100010100    1101001100010101    1101001100010110    1101001100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54035 - 54039

  --1101001100011000    1101001100011001    1101001100011010    1101001100011011    1101001100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54040 - 54044

  --1101001100011101    1101001100011110    1101001100011111    1101001100100000    1101001100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54045 - 54049

  --1101001100100010    1101001100100011    1101001100100100    1101001100100101    1101001100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54050 - 54054

  --1101001100100111    1101001100101000    1101001100101001    1101001100101010    1101001100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54055 - 54059

  --1101001100101100    1101001100101101    1101001100101110    1101001100101111    1101001100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54060 - 54064

  --1101001100110001    1101001100110010    1101001100110011    1101001100110100    1101001100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54065 - 54069

  --1101001100110110    1101001100110111    1101001100111000    1101001100111001    1101001100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54070 - 54074

  --1101001100111011    1101001100111100    1101001100111101    1101001100111110    1101001100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54075 - 54079

  --1101001101000000    1101001101000001    1101001101000010    1101001101000011    1101001101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54080 - 54084

  --1101001101000101    1101001101000110    1101001101000111    1101001101001000    1101001101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54085 - 54089

  --1101001101001010    1101001101001011    1101001101001100    1101001101001101    1101001101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54090 - 54094

  --1101001101001111    1101001101010000    1101001101010001    1101001101010010    1101001101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54095 - 54099

  --1101001101010100    1101001101010101    1101001101010110    1101001101010111    1101001101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54100 - 54104

  --1101001101011001    1101001101011010    1101001101011011    1101001101011100    1101001101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54105 - 54109

  --1101001101011110    1101001101011111    1101001101100000    1101001101100001    1101001101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54110 - 54114

  --1101001101100011    1101001101100100    1101001101100101    1101001101100110    1101001101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54115 - 54119

  --1101001101101000    1101001101101001    1101001101101010    1101001101101011    1101001101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54120 - 54124

  --1101001101101101    1101001101101110    1101001101101111    1101001101110000    1101001101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54125 - 54129

  --1101001101110010    1101001101110011    1101001101110100    1101001101110101    1101001101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54130 - 54134

  --1101001101110111    1101001101111000    1101001101111001    1101001101111010    1101001101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54135 - 54139

  --1101001101111100    1101001101111101    1101001101111110    1101001101111111    1101001110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54140 - 54144

  --1101001110000001    1101001110000010    1101001110000011    1101001110000100    1101001110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54145 - 54149

  --1101001110000110    1101001110000111    1101001110001000    1101001110001001    1101001110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54150 - 54154

  --1101001110001011    1101001110001100    1101001110001101    1101001110001110    1101001110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54155 - 54159

  --1101001110010000    1101001110010001    1101001110010010    1101001110010011    1101001110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54160 - 54164

  --1101001110010101    1101001110010110    1101001110010111    1101001110011000    1101001110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54165 - 54169

  --1101001110011010    1101001110011011    1101001110011100    1101001110011101    1101001110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54170 - 54174

  --1101001110011111    1101001110100000    1101001110100001    1101001110100010    1101001110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54175 - 54179

  --1101001110100100    1101001110100101    1101001110100110    1101001110100111    1101001110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54180 - 54184

  --1101001110101001    1101001110101010    1101001110101011    1101001110101100    1101001110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54185 - 54189

  --1101001110101110    1101001110101111    1101001110110000    1101001110110001    1101001110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54190 - 54194

  --1101001110110011    1101001110110100    1101001110110101    1101001110110110    1101001110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54195 - 54199

  --1101001110111000    1101001110111001    1101001110111010    1101001110111011    1101001110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54200 - 54204

  --1101001110111101    1101001110111110    1101001110111111    1101001111000000    1101001111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54205 - 54209

  --1101001111000010    1101001111000011    1101001111000100    1101001111000101    1101001111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54210 - 54214

  --1101001111000111    1101001111001000    1101001111001001    1101001111001010    1101001111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54215 - 54219

  --1101001111001100    1101001111001101    1101001111001110    1101001111001111    1101001111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54220 - 54224

  --1101001111010001    1101001111010010    1101001111010011    1101001111010100    1101001111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54225 - 54229

  --1101001111010110    1101001111010111    1101001111011000    1101001111011001    1101001111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54230 - 54234

  --1101001111011011    1101001111011100    1101001111011101    1101001111011110    1101001111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54235 - 54239

  --1101001111100000    1101001111100001    1101001111100010    1101001111100011    1101001111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54240 - 54244

  --1101001111100101    1101001111100110    1101001111100111    1101001111101000    1101001111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54245 - 54249

  --1101001111101010    1101001111101011    1101001111101100    1101001111101101    1101001111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54250 - 54254

  --1101001111101111    1101001111110000    1101001111110001    1101001111110010    1101001111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54255 - 54259

  --1101001111110100    1101001111110101    1101001111110110    1101001111110111    1101001111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54260 - 54264

  --1101001111111001    1101001111111010    1101001111111011    1101001111111100    1101001111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54265 - 54269

  --1101001111111110    1101001111111111    1101010000000000    1101010000000001    1101010000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54270 - 54274

  --1101010000000011    1101010000000100    1101010000000101    1101010000000110    1101010000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54275 - 54279

  --1101010000001000    1101010000001001    1101010000001010    1101010000001011    1101010000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54280 - 54284

  --1101010000001101    1101010000001110    1101010000001111    1101010000010000    1101010000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54285 - 54289

  --1101010000010010    1101010000010011    1101010000010100    1101010000010101    1101010000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54290 - 54294

  --1101010000010111    1101010000011000    1101010000011001    1101010000011010    1101010000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54295 - 54299

  --1101010000011100    1101010000011101    1101010000011110    1101010000011111    1101010000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54300 - 54304

  --1101010000100001    1101010000100010    1101010000100011    1101010000100100    1101010000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54305 - 54309

  --1101010000100110    1101010000100111    1101010000101000    1101010000101001    1101010000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54310 - 54314

  --1101010000101011    1101010000101100    1101010000101101    1101010000101110    1101010000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54315 - 54319

  --1101010000110000    1101010000110001    1101010000110010    1101010000110011    1101010000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54320 - 54324

  --1101010000110101    1101010000110110    1101010000110111    1101010000111000    1101010000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54325 - 54329

  --1101010000111010    1101010000111011    1101010000111100    1101010000111101    1101010000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54330 - 54334

  --1101010000111111    1101010001000000    1101010001000001    1101010001000010    1101010001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54335 - 54339

  --1101010001000100    1101010001000101    1101010001000110    1101010001000111    1101010001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54340 - 54344

  --1101010001001001    1101010001001010    1101010001001011    1101010001001100    1101010001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54345 - 54349

  --1101010001001110    1101010001001111    1101010001010000    1101010001010001    1101010001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54350 - 54354

  --1101010001010011    1101010001010100    1101010001010101    1101010001010110    1101010001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54355 - 54359

  --1101010001011000    1101010001011001    1101010001011010    1101010001011011    1101010001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54360 - 54364

  --1101010001011101    1101010001011110    1101010001011111    1101010001100000    1101010001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54365 - 54369

  --1101010001100010    1101010001100011    1101010001100100    1101010001100101    1101010001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54370 - 54374

  --1101010001100111    1101010001101000    1101010001101001    1101010001101010    1101010001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54375 - 54379

  --1101010001101100    1101010001101101    1101010001101110    1101010001101111    1101010001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54380 - 54384

  --1101010001110001    1101010001110010    1101010001110011    1101010001110100    1101010001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54385 - 54389

  --1101010001110110    1101010001110111    1101010001111000    1101010001111001    1101010001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54390 - 54394

  --1101010001111011    1101010001111100    1101010001111101    1101010001111110    1101010001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54395 - 54399

  --1101010010000000    1101010010000001    1101010010000010    1101010010000011    1101010010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54400 - 54404

  --1101010010000101    1101010010000110    1101010010000111    1101010010001000    1101010010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54405 - 54409

  --1101010010001010    1101010010001011    1101010010001100    1101010010001101    1101010010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54410 - 54414

  --1101010010001111    1101010010010000    1101010010010001    1101010010010010    1101010010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54415 - 54419

  --1101010010010100    1101010010010101    1101010010010110    1101010010010111    1101010010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54420 - 54424

  --1101010010011001    1101010010011010    1101010010011011    1101010010011100    1101010010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54425 - 54429

  --1101010010011110    1101010010011111    1101010010100000    1101010010100001    1101010010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54430 - 54434

  --1101010010100011    1101010010100100    1101010010100101    1101010010100110    1101010010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54435 - 54439

  --1101010010101000    1101010010101001    1101010010101010    1101010010101011    1101010010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54440 - 54444

  --1101010010101101    1101010010101110    1101010010101111    1101010010110000    1101010010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54445 - 54449

  --1101010010110010    1101010010110011    1101010010110100    1101010010110101    1101010010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54450 - 54454

  --1101010010110111    1101010010111000    1101010010111001    1101010010111010    1101010010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54455 - 54459

  --1101010010111100    1101010010111101    1101010010111110    1101010010111111    1101010011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54460 - 54464

  --1101010011000001    1101010011000010    1101010011000011    1101010011000100    1101010011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54465 - 54469

  --1101010011000110    1101010011000111    1101010011001000    1101010011001001    1101010011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54470 - 54474

  --1101010011001011    1101010011001100    1101010011001101    1101010011001110    1101010011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54475 - 54479

  --1101010011010000    1101010011010001    1101010011010010    1101010011010011    1101010011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54480 - 54484

  --1101010011010101    1101010011010110    1101010011010111    1101010011011000    1101010011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54485 - 54489

  --1101010011011010    1101010011011011    1101010011011100    1101010011011101    1101010011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54490 - 54494

  --1101010011011111    1101010011100000    1101010011100001    1101010011100010    1101010011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54495 - 54499

  --1101010011100100    1101010011100101    1101010011100110    1101010011100111    1101010011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54500 - 54504

  --1101010011101001    1101010011101010    1101010011101011    1101010011101100    1101010011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54505 - 54509

  --1101010011101110    1101010011101111    1101010011110000    1101010011110001    1101010011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54510 - 54514

  --1101010011110011    1101010011110100    1101010011110101    1101010011110110    1101010011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54515 - 54519

  --1101010011111000    1101010011111001    1101010011111010    1101010011111011    1101010011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54520 - 54524

  --1101010011111101    1101010011111110    1101010011111111    1101010100000000    1101010100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54525 - 54529

  --1101010100000010    1101010100000011    1101010100000100    1101010100000101    1101010100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54530 - 54534

  --1101010100000111    1101010100001000    1101010100001001    1101010100001010    1101010100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54535 - 54539

  --1101010100001100    1101010100001101    1101010100001110    1101010100001111    1101010100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54540 - 54544

  --1101010100010001    1101010100010010    1101010100010011    1101010100010100    1101010100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54545 - 54549

  --1101010100010110    1101010100010111    1101010100011000    1101010100011001    1101010100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54550 - 54554

  --1101010100011011    1101010100011100    1101010100011101    1101010100011110    1101010100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54555 - 54559

  --1101010100100000    1101010100100001    1101010100100010    1101010100100011    1101010100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54560 - 54564

  --1101010100100101    1101010100100110    1101010100100111    1101010100101000    1101010100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54565 - 54569

  --1101010100101010    1101010100101011    1101010100101100    1101010100101101    1101010100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54570 - 54574

  --1101010100101111    1101010100110000    1101010100110001    1101010100110010    1101010100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54575 - 54579

  --1101010100110100    1101010100110101    1101010100110110    1101010100110111    1101010100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54580 - 54584

  --1101010100111001    1101010100111010    1101010100111011    1101010100111100    1101010100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54585 - 54589

  --1101010100111110    1101010100111111    1101010101000000    1101010101000001    1101010101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54590 - 54594

  --1101010101000011    1101010101000100    1101010101000101    1101010101000110    1101010101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54595 - 54599

  --1101010101001000    1101010101001001    1101010101001010    1101010101001011    1101010101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54600 - 54604

  --1101010101001101    1101010101001110    1101010101001111    1101010101010000    1101010101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54605 - 54609

  --1101010101010010    1101010101010011    1101010101010100    1101010101010101    1101010101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54610 - 54614

  --1101010101010111    1101010101011000    1101010101011001    1101010101011010    1101010101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54615 - 54619

  --1101010101011100    1101010101011101    1101010101011110    1101010101011111    1101010101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54620 - 54624

  --1101010101100001    1101010101100010    1101010101100011    1101010101100100    1101010101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54625 - 54629

  --1101010101100110    1101010101100111    1101010101101000    1101010101101001    1101010101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54630 - 54634

  --1101010101101011    1101010101101100    1101010101101101    1101010101101110    1101010101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54635 - 54639

  --1101010101110000    1101010101110001    1101010101110010    1101010101110011    1101010101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54640 - 54644

  --1101010101110101    1101010101110110    1101010101110111    1101010101111000    1101010101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54645 - 54649

  --1101010101111010    1101010101111011    1101010101111100    1101010101111101    1101010101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54650 - 54654

  --1101010101111111    1101010110000000    1101010110000001    1101010110000010    1101010110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54655 - 54659

  --1101010110000100    1101010110000101    1101010110000110    1101010110000111    1101010110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54660 - 54664

  --1101010110001001    1101010110001010    1101010110001011    1101010110001100    1101010110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54665 - 54669

  --1101010110001110    1101010110001111    1101010110010000    1101010110010001    1101010110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54670 - 54674

  --1101010110010011    1101010110010100    1101010110010101    1101010110010110    1101010110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54675 - 54679

  --1101010110011000    1101010110011001    1101010110011010    1101010110011011    1101010110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54680 - 54684

  --1101010110011101    1101010110011110    1101010110011111    1101010110100000    1101010110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54685 - 54689

  --1101010110100010    1101010110100011    1101010110100100    1101010110100101    1101010110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54690 - 54694

  --1101010110100111    1101010110101000    1101010110101001    1101010110101010    1101010110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54695 - 54699

  --1101010110101100    1101010110101101    1101010110101110    1101010110101111    1101010110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54700 - 54704

  --1101010110110001    1101010110110010    1101010110110011    1101010110110100    1101010110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54705 - 54709

  --1101010110110110    1101010110110111    1101010110111000    1101010110111001    1101010110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54710 - 54714

  --1101010110111011    1101010110111100    1101010110111101    1101010110111110    1101010110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54715 - 54719

  --1101010111000000    1101010111000001    1101010111000010    1101010111000011    1101010111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54720 - 54724

  --1101010111000101    1101010111000110    1101010111000111    1101010111001000    1101010111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54725 - 54729

  --1101010111001010    1101010111001011    1101010111001100    1101010111001101    1101010111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54730 - 54734

  --1101010111001111    1101010111010000    1101010111010001    1101010111010010    1101010111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54735 - 54739

  --1101010111010100    1101010111010101    1101010111010110    1101010111010111    1101010111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54740 - 54744

  --1101010111011001    1101010111011010    1101010111011011    1101010111011100    1101010111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54745 - 54749

  --1101010111011110    1101010111011111    1101010111100000    1101010111100001    1101010111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54750 - 54754

  --1101010111100011    1101010111100100    1101010111100101    1101010111100110    1101010111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54755 - 54759

  --1101010111101000    1101010111101001    1101010111101010    1101010111101011    1101010111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54760 - 54764

  --1101010111101101    1101010111101110    1101010111101111    1101010111110000    1101010111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54765 - 54769

  --1101010111110010    1101010111110011    1101010111110100    1101010111110101    1101010111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54770 - 54774

  --1101010111110111    1101010111111000    1101010111111001    1101010111111010    1101010111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54775 - 54779

  --1101010111111100    1101010111111101    1101010111111110    1101010111111111    1101011000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54780 - 54784

  --1101011000000001    1101011000000010    1101011000000011    1101011000000100    1101011000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54785 - 54789

  --1101011000000110    1101011000000111    1101011000001000    1101011000001001    1101011000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54790 - 54794

  --1101011000001011    1101011000001100    1101011000001101    1101011000001110    1101011000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54795 - 54799

  --1101011000010000    1101011000010001    1101011000010010    1101011000010011    1101011000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54800 - 54804

  --1101011000010101    1101011000010110    1101011000010111    1101011000011000    1101011000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54805 - 54809

  --1101011000011010    1101011000011011    1101011000011100    1101011000011101    1101011000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54810 - 54814

  --1101011000011111    1101011000100000    1101011000100001    1101011000100010    1101011000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54815 - 54819

  --1101011000100100    1101011000100101    1101011000100110    1101011000100111    1101011000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54820 - 54824

  --1101011000101001    1101011000101010    1101011000101011    1101011000101100    1101011000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54825 - 54829

  --1101011000101110    1101011000101111    1101011000110000    1101011000110001    1101011000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54830 - 54834

  --1101011000110011    1101011000110100    1101011000110101    1101011000110110    1101011000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54835 - 54839

  --1101011000111000    1101011000111001    1101011000111010    1101011000111011    1101011000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54840 - 54844

  --1101011000111101    1101011000111110    1101011000111111    1101011001000000    1101011001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54845 - 54849

  --1101011001000010    1101011001000011    1101011001000100    1101011001000101    1101011001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54850 - 54854

  --1101011001000111    1101011001001000    1101011001001001    1101011001001010    1101011001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54855 - 54859

  --1101011001001100    1101011001001101    1101011001001110    1101011001001111    1101011001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54860 - 54864

  --1101011001010001    1101011001010010    1101011001010011    1101011001010100    1101011001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54865 - 54869

  --1101011001010110    1101011001010111    1101011001011000    1101011001011001    1101011001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54870 - 54874

  --1101011001011011    1101011001011100    1101011001011101    1101011001011110    1101011001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54875 - 54879

  --1101011001100000    1101011001100001    1101011001100010    1101011001100011    1101011001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54880 - 54884

  --1101011001100101    1101011001100110    1101011001100111    1101011001101000    1101011001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54885 - 54889

  --1101011001101010    1101011001101011    1101011001101100    1101011001101101    1101011001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54890 - 54894

  --1101011001101111    1101011001110000    1101011001110001    1101011001110010    1101011001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54895 - 54899

  --1101011001110100    1101011001110101    1101011001110110    1101011001110111    1101011001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54900 - 54904

  --1101011001111001    1101011001111010    1101011001111011    1101011001111100    1101011001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54905 - 54909

  --1101011001111110    1101011001111111    1101011010000000    1101011010000001    1101011010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54910 - 54914

  --1101011010000011    1101011010000100    1101011010000101    1101011010000110    1101011010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54915 - 54919

  --1101011010001000    1101011010001001    1101011010001010    1101011010001011    1101011010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54920 - 54924

  --1101011010001101    1101011010001110    1101011010001111    1101011010010000    1101011010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54925 - 54929

  --1101011010010010    1101011010010011    1101011010010100    1101011010010101    1101011010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54930 - 54934

  --1101011010010111    1101011010011000    1101011010011001    1101011010011010    1101011010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54935 - 54939

  --1101011010011100    1101011010011101    1101011010011110    1101011010011111    1101011010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54940 - 54944

  --1101011010100001    1101011010100010    1101011010100011    1101011010100100    1101011010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54945 - 54949

  --1101011010100110    1101011010100111    1101011010101000    1101011010101001    1101011010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54950 - 54954

  --1101011010101011    1101011010101100    1101011010101101    1101011010101110    1101011010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54955 - 54959

  --1101011010110000    1101011010110001    1101011010110010    1101011010110011    1101011010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54960 - 54964

  --1101011010110101    1101011010110110    1101011010110111    1101011010111000    1101011010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54965 - 54969

  --1101011010111010    1101011010111011    1101011010111100    1101011010111101    1101011010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54970 - 54974

  --1101011010111111    1101011011000000    1101011011000001    1101011011000010    1101011011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54975 - 54979

  --1101011011000100    1101011011000101    1101011011000110    1101011011000111    1101011011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54980 - 54984

  --1101011011001001    1101011011001010    1101011011001011    1101011011001100    1101011011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54985 - 54989

  --1101011011001110    1101011011001111    1101011011010000    1101011011010001    1101011011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54990 - 54994

  --1101011011010011    1101011011010100    1101011011010101    1101011011010110    1101011011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 54995 - 54999

  --1101011011011000    1101011011011001    1101011011011010    1101011011011011    1101011011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55000 - 55004

  --1101011011011101    1101011011011110    1101011011011111    1101011011100000    1101011011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55005 - 55009

  --1101011011100010    1101011011100011    1101011011100100    1101011011100101    1101011011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55010 - 55014

  --1101011011100111    1101011011101000    1101011011101001    1101011011101010    1101011011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55015 - 55019

  --1101011011101100    1101011011101101    1101011011101110    1101011011101111    1101011011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55020 - 55024

  --1101011011110001    1101011011110010    1101011011110011    1101011011110100    1101011011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55025 - 55029

  --1101011011110110    1101011011110111    1101011011111000    1101011011111001    1101011011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55030 - 55034

  --1101011011111011    1101011011111100    1101011011111101    1101011011111110    1101011011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55035 - 55039

  --1101011100000000    1101011100000001    1101011100000010    1101011100000011    1101011100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55040 - 55044

  --1101011100000101    1101011100000110    1101011100000111    1101011100001000    1101011100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55045 - 55049

  --1101011100001010    1101011100001011    1101011100001100    1101011100001101    1101011100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55050 - 55054

  --1101011100001111    1101011100010000    1101011100010001    1101011100010010    1101011100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55055 - 55059

  --1101011100010100    1101011100010101    1101011100010110    1101011100010111    1101011100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55060 - 55064

  --1101011100011001    1101011100011010    1101011100011011    1101011100011100    1101011100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55065 - 55069

  --1101011100011110    1101011100011111    1101011100100000    1101011100100001    1101011100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55070 - 55074

  --1101011100100011    1101011100100100    1101011100100101    1101011100100110    1101011100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55075 - 55079

  --1101011100101000    1101011100101001    1101011100101010    1101011100101011    1101011100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55080 - 55084

  --1101011100101101    1101011100101110    1101011100101111    1101011100110000    1101011100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55085 - 55089

  --1101011100110010    1101011100110011    1101011100110100    1101011100110101    1101011100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55090 - 55094

  --1101011100110111    1101011100111000    1101011100111001    1101011100111010    1101011100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55095 - 55099

  --1101011100111100    1101011100111101    1101011100111110    1101011100111111    1101011101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55100 - 55104

  --1101011101000001    1101011101000010    1101011101000011    1101011101000100    1101011101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55105 - 55109

  --1101011101000110    1101011101000111    1101011101001000    1101011101001001    1101011101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55110 - 55114

  --1101011101001011    1101011101001100    1101011101001101    1101011101001110    1101011101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55115 - 55119

  --1101011101010000    1101011101010001    1101011101010010    1101011101010011    1101011101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55120 - 55124

  --1101011101010101    1101011101010110    1101011101010111    1101011101011000    1101011101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55125 - 55129

  --1101011101011010    1101011101011011    1101011101011100    1101011101011101    1101011101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55130 - 55134

  --1101011101011111    1101011101100000    1101011101100001    1101011101100010    1101011101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55135 - 55139

  --1101011101100100    1101011101100101    1101011101100110    1101011101100111    1101011101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55140 - 55144

  --1101011101101001    1101011101101010    1101011101101011    1101011101101100    1101011101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55145 - 55149

  --1101011101101110    1101011101101111    1101011101110000    1101011101110001    1101011101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55150 - 55154

  --1101011101110011    1101011101110100    1101011101110101    1101011101110110    1101011101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55155 - 55159

  --1101011101111000    1101011101111001    1101011101111010    1101011101111011    1101011101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55160 - 55164

  --1101011101111101    1101011101111110    1101011101111111    1101011110000000    1101011110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55165 - 55169

  --1101011110000010    1101011110000011    1101011110000100    1101011110000101    1101011110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55170 - 55174

  --1101011110000111    1101011110001000    1101011110001001    1101011110001010    1101011110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55175 - 55179

  --1101011110001100    1101011110001101    1101011110001110    1101011110001111    1101011110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55180 - 55184

  --1101011110010001    1101011110010010    1101011110010011    1101011110010100    1101011110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55185 - 55189

  --1101011110010110    1101011110010111    1101011110011000    1101011110011001    1101011110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55190 - 55194

  --1101011110011011    1101011110011100    1101011110011101    1101011110011110    1101011110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55195 - 55199

  --1101011110100000    1101011110100001    1101011110100010    1101011110100011    1101011110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55200 - 55204

  --1101011110100101    1101011110100110    1101011110100111    1101011110101000    1101011110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55205 - 55209

  --1101011110101010    1101011110101011    1101011110101100    1101011110101101    1101011110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55210 - 55214

  --1101011110101111    1101011110110000    1101011110110001    1101011110110010    1101011110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55215 - 55219

  --1101011110110100    1101011110110101    1101011110110110    1101011110110111    1101011110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55220 - 55224

  --1101011110111001    1101011110111010    1101011110111011    1101011110111100    1101011110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55225 - 55229

  --1101011110111110    1101011110111111    1101011111000000    1101011111000001    1101011111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55230 - 55234

  --1101011111000011    1101011111000100    1101011111000101    1101011111000110    1101011111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55235 - 55239

  --1101011111001000    1101011111001001    1101011111001010    1101011111001011    1101011111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55240 - 55244

  --1101011111001101    1101011111001110    1101011111001111    1101011111010000    1101011111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55245 - 55249

  --1101011111010010    1101011111010011    1101011111010100    1101011111010101    1101011111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55250 - 55254

  --1101011111010111    1101011111011000    1101011111011001    1101011111011010    1101011111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55255 - 55259

  --1101011111011100    1101011111011101    1101011111011110    1101011111011111    1101011111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55260 - 55264

  --1101011111100001    1101011111100010    1101011111100011    1101011111100100    1101011111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55265 - 55269

  --1101011111100110    1101011111100111    1101011111101000    1101011111101001    1101011111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55270 - 55274

  --1101011111101011    1101011111101100    1101011111101101    1101011111101110    1101011111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55275 - 55279

  --1101011111110000    1101011111110001    1101011111110010    1101011111110011    1101011111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55280 - 55284

  --1101011111110101    1101011111110110    1101011111110111    1101011111111000    1101011111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55285 - 55289

  --1101011111111010    1101011111111011    1101011111111100    1101011111111101    1101011111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55290 - 55294

  --1101011111111111    1101100000000000    1101100000000001    1101100000000010    1101100000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55295 - 55299

  --1101100000000100    1101100000000101    1101100000000110    1101100000000111    1101100000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55300 - 55304

  --1101100000001001    1101100000001010    1101100000001011    1101100000001100    1101100000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55305 - 55309

  --1101100000001110    1101100000001111    1101100000010000    1101100000010001    1101100000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55310 - 55314

  --1101100000010011    1101100000010100    1101100000010101    1101100000010110    1101100000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55315 - 55319

  --1101100000011000    1101100000011001    1101100000011010    1101100000011011    1101100000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55320 - 55324

  --1101100000011101    1101100000011110    1101100000011111    1101100000100000    1101100000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55325 - 55329

  --1101100000100010    1101100000100011    1101100000100100    1101100000100101    1101100000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55330 - 55334

  --1101100000100111    1101100000101000    1101100000101001    1101100000101010    1101100000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55335 - 55339

  --1101100000101100    1101100000101101    1101100000101110    1101100000101111    1101100000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55340 - 55344

  --1101100000110001    1101100000110010    1101100000110011    1101100000110100    1101100000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55345 - 55349

  --1101100000110110    1101100000110111    1101100000111000    1101100000111001    1101100000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55350 - 55354

  --1101100000111011    1101100000111100    1101100000111101    1101100000111110    1101100000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55355 - 55359

  --1101100001000000    1101100001000001    1101100001000010    1101100001000011    1101100001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55360 - 55364

  --1101100001000101    1101100001000110    1101100001000111    1101100001001000    1101100001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55365 - 55369

  --1101100001001010    1101100001001011    1101100001001100    1101100001001101    1101100001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55370 - 55374

  --1101100001001111    1101100001010000    1101100001010001    1101100001010010    1101100001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55375 - 55379

  --1101100001010100    1101100001010101    1101100001010110    1101100001010111    1101100001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55380 - 55384

  --1101100001011001    1101100001011010    1101100001011011    1101100001011100    1101100001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55385 - 55389

  --1101100001011110    1101100001011111    1101100001100000    1101100001100001    1101100001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55390 - 55394

  --1101100001100011    1101100001100100    1101100001100101    1101100001100110    1101100001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55395 - 55399

  --1101100001101000    1101100001101001    1101100001101010    1101100001101011    1101100001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55400 - 55404

  --1101100001101101    1101100001101110    1101100001101111    1101100001110000    1101100001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55405 - 55409

  --1101100001110010    1101100001110011    1101100001110100    1101100001110101    1101100001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55410 - 55414

  --1101100001110111    1101100001111000    1101100001111001    1101100001111010    1101100001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55415 - 55419

  --1101100001111100    1101100001111101    1101100001111110    1101100001111111    1101100010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55420 - 55424

  --1101100010000001    1101100010000010    1101100010000011    1101100010000100    1101100010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55425 - 55429

  --1101100010000110    1101100010000111    1101100010001000    1101100010001001    1101100010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55430 - 55434

  --1101100010001011    1101100010001100    1101100010001101    1101100010001110    1101100010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55435 - 55439

  --1101100010010000    1101100010010001    1101100010010010    1101100010010011    1101100010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55440 - 55444

  --1101100010010101    1101100010010110    1101100010010111    1101100010011000    1101100010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55445 - 55449

  --1101100010011010    1101100010011011    1101100010011100    1101100010011101    1101100010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55450 - 55454

  --1101100010011111    1101100010100000    1101100010100001    1101100010100010    1101100010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55455 - 55459

  --1101100010100100    1101100010100101    1101100010100110    1101100010100111    1101100010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55460 - 55464

  --1101100010101001    1101100010101010    1101100010101011    1101100010101100    1101100010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55465 - 55469

  --1101100010101110    1101100010101111    1101100010110000    1101100010110001    1101100010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55470 - 55474

  --1101100010110011    1101100010110100    1101100010110101    1101100010110110    1101100010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55475 - 55479

  --1101100010111000    1101100010111001    1101100010111010    1101100010111011    1101100010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55480 - 55484

  --1101100010111101    1101100010111110    1101100010111111    1101100011000000    1101100011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55485 - 55489

  --1101100011000010    1101100011000011    1101100011000100    1101100011000101    1101100011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55490 - 55494

  --1101100011000111    1101100011001000    1101100011001001    1101100011001010    1101100011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55495 - 55499

  --1101100011001100    1101100011001101    1101100011001110    1101100011001111    1101100011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55500 - 55504

  --1101100011010001    1101100011010010    1101100011010011    1101100011010100    1101100011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55505 - 55509

  --1101100011010110    1101100011010111    1101100011011000    1101100011011001    1101100011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55510 - 55514

  --1101100011011011    1101100011011100    1101100011011101    1101100011011110    1101100011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55515 - 55519

  --1101100011100000    1101100011100001    1101100011100010    1101100011100011    1101100011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55520 - 55524

  --1101100011100101    1101100011100110    1101100011100111    1101100011101000    1101100011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55525 - 55529

  --1101100011101010    1101100011101011    1101100011101100    1101100011101101    1101100011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55530 - 55534

  --1101100011101111    1101100011110000    1101100011110001    1101100011110010    1101100011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55535 - 55539

  --1101100011110100    1101100011110101    1101100011110110    1101100011110111    1101100011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55540 - 55544

  --1101100011111001    1101100011111010    1101100011111011    1101100011111100    1101100011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55545 - 55549

  --1101100011111110    1101100011111111    1101100100000000    1101100100000001    1101100100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55550 - 55554

  --1101100100000011    1101100100000100    1101100100000101    1101100100000110    1101100100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55555 - 55559

  --1101100100001000    1101100100001001    1101100100001010    1101100100001011    1101100100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55560 - 55564

  --1101100100001101    1101100100001110    1101100100001111    1101100100010000    1101100100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55565 - 55569

  --1101100100010010    1101100100010011    1101100100010100    1101100100010101    1101100100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55570 - 55574

  --1101100100010111    1101100100011000    1101100100011001    1101100100011010    1101100100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55575 - 55579

  --1101100100011100    1101100100011101    1101100100011110    1101100100011111    1101100100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55580 - 55584

  --1101100100100001    1101100100100010    1101100100100011    1101100100100100    1101100100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55585 - 55589

  --1101100100100110    1101100100100111    1101100100101000    1101100100101001    1101100100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55590 - 55594

  --1101100100101011    1101100100101100    1101100100101101    1101100100101110    1101100100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55595 - 55599

  --1101100100110000    1101100100110001    1101100100110010    1101100100110011    1101100100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55600 - 55604

  --1101100100110101    1101100100110110    1101100100110111    1101100100111000    1101100100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55605 - 55609

  --1101100100111010    1101100100111011    1101100100111100    1101100100111101    1101100100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55610 - 55614

  --1101100100111111    1101100101000000    1101100101000001    1101100101000010    1101100101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55615 - 55619

  --1101100101000100    1101100101000101    1101100101000110    1101100101000111    1101100101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55620 - 55624

  --1101100101001001    1101100101001010    1101100101001011    1101100101001100    1101100101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55625 - 55629

  --1101100101001110    1101100101001111    1101100101010000    1101100101010001    1101100101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55630 - 55634

  --1101100101010011    1101100101010100    1101100101010101    1101100101010110    1101100101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55635 - 55639

  --1101100101011000    1101100101011001    1101100101011010    1101100101011011    1101100101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55640 - 55644

  --1101100101011101    1101100101011110    1101100101011111    1101100101100000    1101100101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55645 - 55649

  --1101100101100010    1101100101100011    1101100101100100    1101100101100101    1101100101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55650 - 55654

  --1101100101100111    1101100101101000    1101100101101001    1101100101101010    1101100101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55655 - 55659

  --1101100101101100    1101100101101101    1101100101101110    1101100101101111    1101100101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55660 - 55664

  --1101100101110001    1101100101110010    1101100101110011    1101100101110100    1101100101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55665 - 55669

  --1101100101110110    1101100101110111    1101100101111000    1101100101111001    1101100101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55670 - 55674

  --1101100101111011    1101100101111100    1101100101111101    1101100101111110    1101100101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55675 - 55679

  --1101100110000000    1101100110000001    1101100110000010    1101100110000011    1101100110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55680 - 55684

  --1101100110000101    1101100110000110    1101100110000111    1101100110001000    1101100110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55685 - 55689

  --1101100110001010    1101100110001011    1101100110001100    1101100110001101    1101100110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55690 - 55694

  --1101100110001111    1101100110010000    1101100110010001    1101100110010010    1101100110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55695 - 55699

  --1101100110010100    1101100110010101    1101100110010110    1101100110010111    1101100110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55700 - 55704

  --1101100110011001    1101100110011010    1101100110011011    1101100110011100    1101100110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55705 - 55709

  --1101100110011110    1101100110011111    1101100110100000    1101100110100001    1101100110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55710 - 55714

  --1101100110100011    1101100110100100    1101100110100101    1101100110100110    1101100110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55715 - 55719

  --1101100110101000    1101100110101001    1101100110101010    1101100110101011    1101100110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55720 - 55724

  --1101100110101101    1101100110101110    1101100110101111    1101100110110000    1101100110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55725 - 55729

  --1101100110110010    1101100110110011    1101100110110100    1101100110110101    1101100110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55730 - 55734

  --1101100110110111    1101100110111000    1101100110111001    1101100110111010    1101100110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55735 - 55739

  --1101100110111100    1101100110111101    1101100110111110    1101100110111111    1101100111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55740 - 55744

  --1101100111000001    1101100111000010    1101100111000011    1101100111000100    1101100111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55745 - 55749

  --1101100111000110    1101100111000111    1101100111001000    1101100111001001    1101100111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55750 - 55754

  --1101100111001011    1101100111001100    1101100111001101    1101100111001110    1101100111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55755 - 55759

  --1101100111010000    1101100111010001    1101100111010010    1101100111010011    1101100111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55760 - 55764

  --1101100111010101    1101100111010110    1101100111010111    1101100111011000    1101100111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55765 - 55769

  --1101100111011010    1101100111011011    1101100111011100    1101100111011101    1101100111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55770 - 55774

  --1101100111011111    1101100111100000    1101100111100001    1101100111100010    1101100111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55775 - 55779

  --1101100111100100    1101100111100101    1101100111100110    1101100111100111    1101100111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55780 - 55784

  --1101100111101001    1101100111101010    1101100111101011    1101100111101100    1101100111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55785 - 55789

  --1101100111101110    1101100111101111    1101100111110000    1101100111110001    1101100111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55790 - 55794

  --1101100111110011    1101100111110100    1101100111110101    1101100111110110    1101100111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55795 - 55799

  --1101100111111000    1101100111111001    1101100111111010    1101100111111011    1101100111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55800 - 55804

  --1101100111111101    1101100111111110    1101100111111111    1101101000000000    1101101000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55805 - 55809

  --1101101000000010    1101101000000011    1101101000000100    1101101000000101    1101101000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55810 - 55814

  --1101101000000111    1101101000001000    1101101000001001    1101101000001010    1101101000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55815 - 55819

  --1101101000001100    1101101000001101    1101101000001110    1101101000001111    1101101000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55820 - 55824

  --1101101000010001    1101101000010010    1101101000010011    1101101000010100    1101101000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55825 - 55829

  --1101101000010110    1101101000010111    1101101000011000    1101101000011001    1101101000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55830 - 55834

  --1101101000011011    1101101000011100    1101101000011101    1101101000011110    1101101000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55835 - 55839

  --1101101000100000    1101101000100001    1101101000100010    1101101000100011    1101101000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55840 - 55844

  --1101101000100101    1101101000100110    1101101000100111    1101101000101000    1101101000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55845 - 55849

  --1101101000101010    1101101000101011    1101101000101100    1101101000101101    1101101000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55850 - 55854

  --1101101000101111    1101101000110000    1101101000110001    1101101000110010    1101101000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55855 - 55859

  --1101101000110100    1101101000110101    1101101000110110    1101101000110111    1101101000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55860 - 55864

  --1101101000111001    1101101000111010    1101101000111011    1101101000111100    1101101000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55865 - 55869

  --1101101000111110    1101101000111111    1101101001000000    1101101001000001    1101101001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55870 - 55874

  --1101101001000011    1101101001000100    1101101001000101    1101101001000110    1101101001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55875 - 55879

  --1101101001001000    1101101001001001    1101101001001010    1101101001001011    1101101001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55880 - 55884

  --1101101001001101    1101101001001110    1101101001001111    1101101001010000    1101101001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55885 - 55889

  --1101101001010010    1101101001010011    1101101001010100    1101101001010101    1101101001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55890 - 55894

  --1101101001010111    1101101001011000    1101101001011001    1101101001011010    1101101001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55895 - 55899

  --1101101001011100    1101101001011101    1101101001011110    1101101001011111    1101101001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55900 - 55904

  --1101101001100001    1101101001100010    1101101001100011    1101101001100100    1101101001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55905 - 55909

  --1101101001100110    1101101001100111    1101101001101000    1101101001101001    1101101001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55910 - 55914

  --1101101001101011    1101101001101100    1101101001101101    1101101001101110    1101101001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55915 - 55919

  --1101101001110000    1101101001110001    1101101001110010    1101101001110011    1101101001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55920 - 55924

  --1101101001110101    1101101001110110    1101101001110111    1101101001111000    1101101001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55925 - 55929

  --1101101001111010    1101101001111011    1101101001111100    1101101001111101    1101101001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55930 - 55934

  --1101101001111111    1101101010000000    1101101010000001    1101101010000010    1101101010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55935 - 55939

  --1101101010000100    1101101010000101    1101101010000110    1101101010000111    1101101010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55940 - 55944

  --1101101010001001    1101101010001010    1101101010001011    1101101010001100    1101101010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55945 - 55949

  --1101101010001110    1101101010001111    1101101010010000    1101101010010001    1101101010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55950 - 55954

  --1101101010010011    1101101010010100    1101101010010101    1101101010010110    1101101010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55955 - 55959

  --1101101010011000    1101101010011001    1101101010011010    1101101010011011    1101101010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55960 - 55964

  --1101101010011101    1101101010011110    1101101010011111    1101101010100000    1101101010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55965 - 55969

  --1101101010100010    1101101010100011    1101101010100100    1101101010100101    1101101010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55970 - 55974

  --1101101010100111    1101101010101000    1101101010101001    1101101010101010    1101101010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55975 - 55979

  --1101101010101100    1101101010101101    1101101010101110    1101101010101111    1101101010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55980 - 55984

  --1101101010110001    1101101010110010    1101101010110011    1101101010110100    1101101010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55985 - 55989

  --1101101010110110    1101101010110111    1101101010111000    1101101010111001    1101101010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55990 - 55994

  --1101101010111011    1101101010111100    1101101010111101    1101101010111110    1101101010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 55995 - 55999

  --1101101011000000    1101101011000001    1101101011000010    1101101011000011    1101101011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56000 - 56004

  --1101101011000101    1101101011000110    1101101011000111    1101101011001000    1101101011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56005 - 56009

  --1101101011001010    1101101011001011    1101101011001100    1101101011001101    1101101011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56010 - 56014

  --1101101011001111    1101101011010000    1101101011010001    1101101011010010    1101101011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56015 - 56019

  --1101101011010100    1101101011010101    1101101011010110    1101101011010111    1101101011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56020 - 56024

  --1101101011011001    1101101011011010    1101101011011011    1101101011011100    1101101011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56025 - 56029

  --1101101011011110    1101101011011111    1101101011100000    1101101011100001    1101101011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56030 - 56034

  --1101101011100011    1101101011100100    1101101011100101    1101101011100110    1101101011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56035 - 56039

  --1101101011101000    1101101011101001    1101101011101010    1101101011101011    1101101011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56040 - 56044

  --1101101011101101    1101101011101110    1101101011101111    1101101011110000    1101101011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56045 - 56049

  --1101101011110010    1101101011110011    1101101011110100    1101101011110101    1101101011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56050 - 56054

  --1101101011110111    1101101011111000    1101101011111001    1101101011111010    1101101011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56055 - 56059

  --1101101011111100    1101101011111101    1101101011111110    1101101011111111    1101101100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56060 - 56064

  --1101101100000001    1101101100000010    1101101100000011    1101101100000100    1101101100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56065 - 56069

  --1101101100000110    1101101100000111    1101101100001000    1101101100001001    1101101100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56070 - 56074

  --1101101100001011    1101101100001100    1101101100001101    1101101100001110    1101101100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56075 - 56079

  --1101101100010000    1101101100010001    1101101100010010    1101101100010011    1101101100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56080 - 56084

  --1101101100010101    1101101100010110    1101101100010111    1101101100011000    1101101100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56085 - 56089

  --1101101100011010    1101101100011011    1101101100011100    1101101100011101    1101101100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56090 - 56094

  --1101101100011111    1101101100100000    1101101100100001    1101101100100010    1101101100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56095 - 56099

  --1101101100100100    1101101100100101    1101101100100110    1101101100100111    1101101100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56100 - 56104

  --1101101100101001    1101101100101010    1101101100101011    1101101100101100    1101101100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56105 - 56109

  --1101101100101110    1101101100101111    1101101100110000    1101101100110001    1101101100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56110 - 56114

  --1101101100110011    1101101100110100    1101101100110101    1101101100110110    1101101100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56115 - 56119

  --1101101100111000    1101101100111001    1101101100111010    1101101100111011    1101101100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56120 - 56124

  --1101101100111101    1101101100111110    1101101100111111    1101101101000000    1101101101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56125 - 56129

  --1101101101000010    1101101101000011    1101101101000100    1101101101000101    1101101101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56130 - 56134

  --1101101101000111    1101101101001000    1101101101001001    1101101101001010    1101101101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56135 - 56139

  --1101101101001100    1101101101001101    1101101101001110    1101101101001111    1101101101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56140 - 56144

  --1101101101010001    1101101101010010    1101101101010011    1101101101010100    1101101101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56145 - 56149

  --1101101101010110    1101101101010111    1101101101011000    1101101101011001    1101101101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56150 - 56154

  --1101101101011011    1101101101011100    1101101101011101    1101101101011110    1101101101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56155 - 56159

  --1101101101100000    1101101101100001    1101101101100010    1101101101100011    1101101101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56160 - 56164

  --1101101101100101    1101101101100110    1101101101100111    1101101101101000    1101101101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56165 - 56169

  --1101101101101010    1101101101101011    1101101101101100    1101101101101101    1101101101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56170 - 56174

  --1101101101101111    1101101101110000    1101101101110001    1101101101110010    1101101101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56175 - 56179

  --1101101101110100    1101101101110101    1101101101110110    1101101101110111    1101101101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56180 - 56184

  --1101101101111001    1101101101111010    1101101101111011    1101101101111100    1101101101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56185 - 56189

  --1101101101111110    1101101101111111    1101101110000000    1101101110000001    1101101110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56190 - 56194

  --1101101110000011    1101101110000100    1101101110000101    1101101110000110    1101101110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56195 - 56199

  --1101101110001000    1101101110001001    1101101110001010    1101101110001011    1101101110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56200 - 56204

  --1101101110001101    1101101110001110    1101101110001111    1101101110010000    1101101110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56205 - 56209

  --1101101110010010    1101101110010011    1101101110010100    1101101110010101    1101101110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56210 - 56214

  --1101101110010111    1101101110011000    1101101110011001    1101101110011010    1101101110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56215 - 56219

  --1101101110011100    1101101110011101    1101101110011110    1101101110011111    1101101110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56220 - 56224

  --1101101110100001    1101101110100010    1101101110100011    1101101110100100    1101101110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56225 - 56229

  --1101101110100110    1101101110100111    1101101110101000    1101101110101001    1101101110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56230 - 56234

  --1101101110101011    1101101110101100    1101101110101101    1101101110101110    1101101110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56235 - 56239

  --1101101110110000    1101101110110001    1101101110110010    1101101110110011    1101101110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56240 - 56244

  --1101101110110101    1101101110110110    1101101110110111    1101101110111000    1101101110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56245 - 56249

  --1101101110111010    1101101110111011    1101101110111100    1101101110111101    1101101110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56250 - 56254

  --1101101110111111    1101101111000000    1101101111000001    1101101111000010    1101101111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56255 - 56259

  --1101101111000100    1101101111000101    1101101111000110    1101101111000111    1101101111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56260 - 56264

  --1101101111001001    1101101111001010    1101101111001011    1101101111001100    1101101111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56265 - 56269

  --1101101111001110    1101101111001111    1101101111010000    1101101111010001    1101101111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56270 - 56274

  --1101101111010011    1101101111010100    1101101111010101    1101101111010110    1101101111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56275 - 56279

  --1101101111011000    1101101111011001    1101101111011010    1101101111011011    1101101111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56280 - 56284

  --1101101111011101    1101101111011110    1101101111011111    1101101111100000    1101101111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56285 - 56289

  --1101101111100010    1101101111100011    1101101111100100    1101101111100101    1101101111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56290 - 56294

  --1101101111100111    1101101111101000    1101101111101001    1101101111101010    1101101111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56295 - 56299

  --1101101111101100    1101101111101101    1101101111101110    1101101111101111    1101101111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56300 - 56304

  --1101101111110001    1101101111110010    1101101111110011    1101101111110100    1101101111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56305 - 56309

  --1101101111110110    1101101111110111    1101101111111000    1101101111111001    1101101111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56310 - 56314

  --1101101111111011    1101101111111100    1101101111111101    1101101111111110    1101101111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56315 - 56319

  --1101110000000000    1101110000000001    1101110000000010    1101110000000011    1101110000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56320 - 56324

  --1101110000000101    1101110000000110    1101110000000111    1101110000001000    1101110000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56325 - 56329

  --1101110000001010    1101110000001011    1101110000001100    1101110000001101    1101110000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56330 - 56334

  --1101110000001111    1101110000010000    1101110000010001    1101110000010010    1101110000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56335 - 56339

  --1101110000010100    1101110000010101    1101110000010110    1101110000010111    1101110000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56340 - 56344

  --1101110000011001    1101110000011010    1101110000011011    1101110000011100    1101110000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56345 - 56349

  --1101110000011110    1101110000011111    1101110000100000    1101110000100001    1101110000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56350 - 56354

  --1101110000100011    1101110000100100    1101110000100101    1101110000100110    1101110000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56355 - 56359

  --1101110000101000    1101110000101001    1101110000101010    1101110000101011    1101110000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56360 - 56364

  --1101110000101101    1101110000101110    1101110000101111    1101110000110000    1101110000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56365 - 56369

  --1101110000110010    1101110000110011    1101110000110100    1101110000110101    1101110000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56370 - 56374

  --1101110000110111    1101110000111000    1101110000111001    1101110000111010    1101110000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56375 - 56379

  --1101110000111100    1101110000111101    1101110000111110    1101110000111111    1101110001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56380 - 56384

  --1101110001000001    1101110001000010    1101110001000011    1101110001000100    1101110001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56385 - 56389

  --1101110001000110    1101110001000111    1101110001001000    1101110001001001    1101110001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56390 - 56394

  --1101110001001011    1101110001001100    1101110001001101    1101110001001110    1101110001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56395 - 56399

  --1101110001010000    1101110001010001    1101110001010010    1101110001010011    1101110001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56400 - 56404

  --1101110001010101    1101110001010110    1101110001010111    1101110001011000    1101110001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56405 - 56409

  --1101110001011010    1101110001011011    1101110001011100    1101110001011101    1101110001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56410 - 56414

  --1101110001011111    1101110001100000    1101110001100001    1101110001100010    1101110001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56415 - 56419

  --1101110001100100    1101110001100101    1101110001100110    1101110001100111    1101110001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56420 - 56424

  --1101110001101001    1101110001101010    1101110001101011    1101110001101100    1101110001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56425 - 56429

  --1101110001101110    1101110001101111    1101110001110000    1101110001110001    1101110001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56430 - 56434

  --1101110001110011    1101110001110100    1101110001110101    1101110001110110    1101110001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56435 - 56439

  --1101110001111000    1101110001111001    1101110001111010    1101110001111011    1101110001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56440 - 56444

  --1101110001111101    1101110001111110    1101110001111111    1101110010000000    1101110010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56445 - 56449

  --1101110010000010    1101110010000011    1101110010000100    1101110010000101    1101110010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56450 - 56454

  --1101110010000111    1101110010001000    1101110010001001    1101110010001010    1101110010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56455 - 56459

  --1101110010001100    1101110010001101    1101110010001110    1101110010001111    1101110010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56460 - 56464

  --1101110010010001    1101110010010010    1101110010010011    1101110010010100    1101110010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56465 - 56469

  --1101110010010110    1101110010010111    1101110010011000    1101110010011001    1101110010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56470 - 56474

  --1101110010011011    1101110010011100    1101110010011101    1101110010011110    1101110010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56475 - 56479

  --1101110010100000    1101110010100001    1101110010100010    1101110010100011    1101110010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56480 - 56484

  --1101110010100101    1101110010100110    1101110010100111    1101110010101000    1101110010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56485 - 56489

  --1101110010101010    1101110010101011    1101110010101100    1101110010101101    1101110010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56490 - 56494

  --1101110010101111    1101110010110000    1101110010110001    1101110010110010    1101110010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56495 - 56499

  --1101110010110100    1101110010110101    1101110010110110    1101110010110111    1101110010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56500 - 56504

  --1101110010111001    1101110010111010    1101110010111011    1101110010111100    1101110010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56505 - 56509

  --1101110010111110    1101110010111111    1101110011000000    1101110011000001    1101110011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56510 - 56514

  --1101110011000011    1101110011000100    1101110011000101    1101110011000110    1101110011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56515 - 56519

  --1101110011001000    1101110011001001    1101110011001010    1101110011001011    1101110011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56520 - 56524

  --1101110011001101    1101110011001110    1101110011001111    1101110011010000    1101110011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56525 - 56529

  --1101110011010010    1101110011010011    1101110011010100    1101110011010101    1101110011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56530 - 56534

  --1101110011010111    1101110011011000    1101110011011001    1101110011011010    1101110011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56535 - 56539

  --1101110011011100    1101110011011101    1101110011011110    1101110011011111    1101110011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56540 - 56544

  --1101110011100001    1101110011100010    1101110011100011    1101110011100100    1101110011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56545 - 56549

  --1101110011100110    1101110011100111    1101110011101000    1101110011101001    1101110011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56550 - 56554

  --1101110011101011    1101110011101100    1101110011101101    1101110011101110    1101110011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56555 - 56559

  --1101110011110000    1101110011110001    1101110011110010    1101110011110011    1101110011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56560 - 56564

  --1101110011110101    1101110011110110    1101110011110111    1101110011111000    1101110011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56565 - 56569

  --1101110011111010    1101110011111011    1101110011111100    1101110011111101    1101110011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56570 - 56574

  --1101110011111111    1101110100000000    1101110100000001    1101110100000010    1101110100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56575 - 56579

  --1101110100000100    1101110100000101    1101110100000110    1101110100000111    1101110100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56580 - 56584

  --1101110100001001    1101110100001010    1101110100001011    1101110100001100    1101110100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56585 - 56589

  --1101110100001110    1101110100001111    1101110100010000    1101110100010001    1101110100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56590 - 56594

  --1101110100010011    1101110100010100    1101110100010101    1101110100010110    1101110100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56595 - 56599

  --1101110100011000    1101110100011001    1101110100011010    1101110100011011    1101110100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56600 - 56604

  --1101110100011101    1101110100011110    1101110100011111    1101110100100000    1101110100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56605 - 56609

  --1101110100100010    1101110100100011    1101110100100100    1101110100100101    1101110100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56610 - 56614

  --1101110100100111    1101110100101000    1101110100101001    1101110100101010    1101110100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56615 - 56619

  --1101110100101100    1101110100101101    1101110100101110    1101110100101111    1101110100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56620 - 56624

  --1101110100110001    1101110100110010    1101110100110011    1101110100110100    1101110100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56625 - 56629

  --1101110100110110    1101110100110111    1101110100111000    1101110100111001    1101110100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56630 - 56634

  --1101110100111011    1101110100111100    1101110100111101    1101110100111110    1101110100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56635 - 56639

  --1101110101000000    1101110101000001    1101110101000010    1101110101000011    1101110101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56640 - 56644

  --1101110101000101    1101110101000110    1101110101000111    1101110101001000    1101110101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56645 - 56649

  --1101110101001010    1101110101001011    1101110101001100    1101110101001101    1101110101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56650 - 56654

  --1101110101001111    1101110101010000    1101110101010001    1101110101010010    1101110101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56655 - 56659

  --1101110101010100    1101110101010101    1101110101010110    1101110101010111    1101110101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56660 - 56664

  --1101110101011001    1101110101011010    1101110101011011    1101110101011100    1101110101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56665 - 56669

  --1101110101011110    1101110101011111    1101110101100000    1101110101100001    1101110101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56670 - 56674

  --1101110101100011    1101110101100100    1101110101100101    1101110101100110    1101110101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56675 - 56679

  --1101110101101000    1101110101101001    1101110101101010    1101110101101011    1101110101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56680 - 56684

  --1101110101101101    1101110101101110    1101110101101111    1101110101110000    1101110101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56685 - 56689

  --1101110101110010    1101110101110011    1101110101110100    1101110101110101    1101110101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56690 - 56694

  --1101110101110111    1101110101111000    1101110101111001    1101110101111010    1101110101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56695 - 56699

  --1101110101111100    1101110101111101    1101110101111110    1101110101111111    1101110110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56700 - 56704

  --1101110110000001    1101110110000010    1101110110000011    1101110110000100    1101110110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56705 - 56709

  --1101110110000110    1101110110000111    1101110110001000    1101110110001001    1101110110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56710 - 56714

  --1101110110001011    1101110110001100    1101110110001101    1101110110001110    1101110110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56715 - 56719

  --1101110110010000    1101110110010001    1101110110010010    1101110110010011    1101110110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56720 - 56724

  --1101110110010101    1101110110010110    1101110110010111    1101110110011000    1101110110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56725 - 56729

  --1101110110011010    1101110110011011    1101110110011100    1101110110011101    1101110110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56730 - 56734

  --1101110110011111    1101110110100000    1101110110100001    1101110110100010    1101110110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56735 - 56739

  --1101110110100100    1101110110100101    1101110110100110    1101110110100111    1101110110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56740 - 56744

  --1101110110101001    1101110110101010    1101110110101011    1101110110101100    1101110110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56745 - 56749

  --1101110110101110    1101110110101111    1101110110110000    1101110110110001    1101110110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56750 - 56754

  --1101110110110011    1101110110110100    1101110110110101    1101110110110110    1101110110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56755 - 56759

  --1101110110111000    1101110110111001    1101110110111010    1101110110111011    1101110110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56760 - 56764

  --1101110110111101    1101110110111110    1101110110111111    1101110111000000    1101110111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56765 - 56769

  --1101110111000010    1101110111000011    1101110111000100    1101110111000101    1101110111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56770 - 56774

  --1101110111000111    1101110111001000    1101110111001001    1101110111001010    1101110111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56775 - 56779

  --1101110111001100    1101110111001101    1101110111001110    1101110111001111    1101110111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56780 - 56784

  --1101110111010001    1101110111010010    1101110111010011    1101110111010100    1101110111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56785 - 56789

  --1101110111010110    1101110111010111    1101110111011000    1101110111011001    1101110111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56790 - 56794

  --1101110111011011    1101110111011100    1101110111011101    1101110111011110    1101110111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56795 - 56799

  --1101110111100000    1101110111100001    1101110111100010    1101110111100011    1101110111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56800 - 56804

  --1101110111100101    1101110111100110    1101110111100111    1101110111101000    1101110111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56805 - 56809

  --1101110111101010    1101110111101011    1101110111101100    1101110111101101    1101110111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56810 - 56814

  --1101110111101111    1101110111110000    1101110111110001    1101110111110010    1101110111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56815 - 56819

  --1101110111110100    1101110111110101    1101110111110110    1101110111110111    1101110111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56820 - 56824

  --1101110111111001    1101110111111010    1101110111111011    1101110111111100    1101110111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56825 - 56829

  --1101110111111110    1101110111111111    1101111000000000    1101111000000001    1101111000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56830 - 56834

  --1101111000000011    1101111000000100    1101111000000101    1101111000000110    1101111000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56835 - 56839

  --1101111000001000    1101111000001001    1101111000001010    1101111000001011    1101111000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56840 - 56844

  --1101111000001101    1101111000001110    1101111000001111    1101111000010000    1101111000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56845 - 56849

  --1101111000010010    1101111000010011    1101111000010100    1101111000010101    1101111000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56850 - 56854

  --1101111000010111    1101111000011000    1101111000011001    1101111000011010    1101111000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56855 - 56859

  --1101111000011100    1101111000011101    1101111000011110    1101111000011111    1101111000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56860 - 56864

  --1101111000100001    1101111000100010    1101111000100011    1101111000100100    1101111000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56865 - 56869

  --1101111000100110    1101111000100111    1101111000101000    1101111000101001    1101111000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56870 - 56874

  --1101111000101011    1101111000101100    1101111000101101    1101111000101110    1101111000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56875 - 56879

  --1101111000110000    1101111000110001    1101111000110010    1101111000110011    1101111000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56880 - 56884

  --1101111000110101    1101111000110110    1101111000110111    1101111000111000    1101111000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56885 - 56889

  --1101111000111010    1101111000111011    1101111000111100    1101111000111101    1101111000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56890 - 56894

  --1101111000111111    1101111001000000    1101111001000001    1101111001000010    1101111001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56895 - 56899

  --1101111001000100    1101111001000101    1101111001000110    1101111001000111    1101111001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56900 - 56904

  --1101111001001001    1101111001001010    1101111001001011    1101111001001100    1101111001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56905 - 56909

  --1101111001001110    1101111001001111    1101111001010000    1101111001010001    1101111001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56910 - 56914

  --1101111001010011    1101111001010100    1101111001010101    1101111001010110    1101111001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56915 - 56919

  --1101111001011000    1101111001011001    1101111001011010    1101111001011011    1101111001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56920 - 56924

  --1101111001011101    1101111001011110    1101111001011111    1101111001100000    1101111001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56925 - 56929

  --1101111001100010    1101111001100011    1101111001100100    1101111001100101    1101111001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56930 - 56934

  --1101111001100111    1101111001101000    1101111001101001    1101111001101010    1101111001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56935 - 56939

  --1101111001101100    1101111001101101    1101111001101110    1101111001101111    1101111001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56940 - 56944

  --1101111001110001    1101111001110010    1101111001110011    1101111001110100    1101111001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56945 - 56949

  --1101111001110110    1101111001110111    1101111001111000    1101111001111001    1101111001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56950 - 56954

  --1101111001111011    1101111001111100    1101111001111101    1101111001111110    1101111001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56955 - 56959

  --1101111010000000    1101111010000001    1101111010000010    1101111010000011    1101111010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56960 - 56964

  --1101111010000101    1101111010000110    1101111010000111    1101111010001000    1101111010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56965 - 56969

  --1101111010001010    1101111010001011    1101111010001100    1101111010001101    1101111010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56970 - 56974

  --1101111010001111    1101111010010000    1101111010010001    1101111010010010    1101111010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56975 - 56979

  --1101111010010100    1101111010010101    1101111010010110    1101111010010111    1101111010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56980 - 56984

  --1101111010011001    1101111010011010    1101111010011011    1101111010011100    1101111010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56985 - 56989

  --1101111010011110    1101111010011111    1101111010100000    1101111010100001    1101111010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56990 - 56994

  --1101111010100011    1101111010100100    1101111010100101    1101111010100110    1101111010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 56995 - 56999

  --1101111010101000    1101111010101001    1101111010101010    1101111010101011    1101111010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57000 - 57004

  --1101111010101101    1101111010101110    1101111010101111    1101111010110000    1101111010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57005 - 57009

  --1101111010110010    1101111010110011    1101111010110100    1101111010110101    1101111010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57010 - 57014

  --1101111010110111    1101111010111000    1101111010111001    1101111010111010    1101111010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57015 - 57019

  --1101111010111100    1101111010111101    1101111010111110    1101111010111111    1101111011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57020 - 57024

  --1101111011000001    1101111011000010    1101111011000011    1101111011000100    1101111011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57025 - 57029

  --1101111011000110    1101111011000111    1101111011001000    1101111011001001    1101111011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57030 - 57034

  --1101111011001011    1101111011001100    1101111011001101    1101111011001110    1101111011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57035 - 57039

  --1101111011010000    1101111011010001    1101111011010010    1101111011010011    1101111011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57040 - 57044

  --1101111011010101    1101111011010110    1101111011010111    1101111011011000    1101111011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57045 - 57049

  --1101111011011010    1101111011011011    1101111011011100    1101111011011101    1101111011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57050 - 57054

  --1101111011011111    1101111011100000    1101111011100001    1101111011100010    1101111011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57055 - 57059

  --1101111011100100    1101111011100101    1101111011100110    1101111011100111    1101111011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57060 - 57064

  --1101111011101001    1101111011101010    1101111011101011    1101111011101100    1101111011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57065 - 57069

  --1101111011101110    1101111011101111    1101111011110000    1101111011110001    1101111011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57070 - 57074

  --1101111011110011    1101111011110100    1101111011110101    1101111011110110    1101111011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57075 - 57079

  --1101111011111000    1101111011111001    1101111011111010    1101111011111011    1101111011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57080 - 57084

  --1101111011111101    1101111011111110    1101111011111111    1101111100000000    1101111100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57085 - 57089

  --1101111100000010    1101111100000011    1101111100000100    1101111100000101    1101111100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57090 - 57094

  --1101111100000111    1101111100001000    1101111100001001    1101111100001010    1101111100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57095 - 57099

  --1101111100001100    1101111100001101    1101111100001110    1101111100001111    1101111100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57100 - 57104

  --1101111100010001    1101111100010010    1101111100010011    1101111100010100    1101111100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57105 - 57109

  --1101111100010110    1101111100010111    1101111100011000    1101111100011001    1101111100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57110 - 57114

  --1101111100011011    1101111100011100    1101111100011101    1101111100011110    1101111100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57115 - 57119

  --1101111100100000    1101111100100001    1101111100100010    1101111100100011    1101111100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57120 - 57124

  --1101111100100101    1101111100100110    1101111100100111    1101111100101000    1101111100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57125 - 57129

  --1101111100101010    1101111100101011    1101111100101100    1101111100101101    1101111100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57130 - 57134

  --1101111100101111    1101111100110000    1101111100110001    1101111100110010    1101111100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57135 - 57139

  --1101111100110100    1101111100110101    1101111100110110    1101111100110111    1101111100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57140 - 57144

  --1101111100111001    1101111100111010    1101111100111011    1101111100111100    1101111100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57145 - 57149

  --1101111100111110    1101111100111111    1101111101000000    1101111101000001    1101111101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57150 - 57154

  --1101111101000011    1101111101000100    1101111101000101    1101111101000110    1101111101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57155 - 57159

  --1101111101001000    1101111101001001    1101111101001010    1101111101001011    1101111101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57160 - 57164

  --1101111101001101    1101111101001110    1101111101001111    1101111101010000    1101111101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57165 - 57169

  --1101111101010010    1101111101010011    1101111101010100    1101111101010101    1101111101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57170 - 57174

  --1101111101010111    1101111101011000    1101111101011001    1101111101011010    1101111101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57175 - 57179

  --1101111101011100    1101111101011101    1101111101011110    1101111101011111    1101111101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57180 - 57184

  --1101111101100001    1101111101100010    1101111101100011    1101111101100100    1101111101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57185 - 57189

  --1101111101100110    1101111101100111    1101111101101000    1101111101101001    1101111101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57190 - 57194

  --1101111101101011    1101111101101100    1101111101101101    1101111101101110    1101111101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57195 - 57199

  --1101111101110000    1101111101110001    1101111101110010    1101111101110011    1101111101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57200 - 57204

  --1101111101110101    1101111101110110    1101111101110111    1101111101111000    1101111101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57205 - 57209

  --1101111101111010    1101111101111011    1101111101111100    1101111101111101    1101111101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57210 - 57214

  --1101111101111111    1101111110000000    1101111110000001    1101111110000010    1101111110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57215 - 57219

  --1101111110000100    1101111110000101    1101111110000110    1101111110000111    1101111110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57220 - 57224

  --1101111110001001    1101111110001010    1101111110001011    1101111110001100    1101111110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57225 - 57229

  --1101111110001110    1101111110001111    1101111110010000    1101111110010001    1101111110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57230 - 57234

  --1101111110010011    1101111110010100    1101111110010101    1101111110010110    1101111110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57235 - 57239

  --1101111110011000    1101111110011001    1101111110011010    1101111110011011    1101111110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57240 - 57244

  --1101111110011101    1101111110011110    1101111110011111    1101111110100000    1101111110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57245 - 57249

  --1101111110100010    1101111110100011    1101111110100100    1101111110100101    1101111110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57250 - 57254

  --1101111110100111    1101111110101000    1101111110101001    1101111110101010    1101111110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57255 - 57259

  --1101111110101100    1101111110101101    1101111110101110    1101111110101111    1101111110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57260 - 57264

  --1101111110110001    1101111110110010    1101111110110011    1101111110110100    1101111110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57265 - 57269

  --1101111110110110    1101111110110111    1101111110111000    1101111110111001    1101111110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57270 - 57274

  --1101111110111011    1101111110111100    1101111110111101    1101111110111110    1101111110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57275 - 57279

  --1101111111000000    1101111111000001    1101111111000010    1101111111000011    1101111111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57280 - 57284

  --1101111111000101    1101111111000110    1101111111000111    1101111111001000    1101111111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57285 - 57289

  --1101111111001010    1101111111001011    1101111111001100    1101111111001101    1101111111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57290 - 57294

  --1101111111001111    1101111111010000    1101111111010001    1101111111010010    1101111111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57295 - 57299

  --1101111111010100    1101111111010101    1101111111010110    1101111111010111    1101111111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57300 - 57304

  --1101111111011001    1101111111011010    1101111111011011    1101111111011100    1101111111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57305 - 57309

  --1101111111011110    1101111111011111    1101111111100000    1101111111100001    1101111111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57310 - 57314

  --1101111111100011    1101111111100100    1101111111100101    1101111111100110    1101111111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57315 - 57319

  --1101111111101000    1101111111101001    1101111111101010    1101111111101011    1101111111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57320 - 57324

  --1101111111101101    1101111111101110    1101111111101111    1101111111110000    1101111111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57325 - 57329

  --1101111111110010    1101111111110011    1101111111110100    1101111111110101    1101111111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57330 - 57334

  --1101111111110111    1101111111111000    1101111111111001    1101111111111010    1101111111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57335 - 57339

  --1101111111111100    1101111111111101    1101111111111110    1101111111111111    1110000000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57340 - 57344

  --1110000000000001    1110000000000010    1110000000000011    1110000000000100    1110000000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57345 - 57349

  --1110000000000110    1110000000000111    1110000000001000    1110000000001001    1110000000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57350 - 57354

  --1110000000001011    1110000000001100    1110000000001101    1110000000001110    1110000000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57355 - 57359

  --1110000000010000    1110000000010001    1110000000010010    1110000000010011    1110000000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57360 - 57364

  --1110000000010101    1110000000010110    1110000000010111    1110000000011000    1110000000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57365 - 57369

  --1110000000011010    1110000000011011    1110000000011100    1110000000011101    1110000000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57370 - 57374

  --1110000000011111    1110000000100000    1110000000100001    1110000000100010    1110000000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57375 - 57379

  --1110000000100100    1110000000100101    1110000000100110    1110000000100111    1110000000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57380 - 57384

  --1110000000101001    1110000000101010    1110000000101011    1110000000101100    1110000000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57385 - 57389

  --1110000000101110    1110000000101111    1110000000110000    1110000000110001    1110000000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57390 - 57394

  --1110000000110011    1110000000110100    1110000000110101    1110000000110110    1110000000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57395 - 57399

  --1110000000111000    1110000000111001    1110000000111010    1110000000111011    1110000000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57400 - 57404

  --1110000000111101    1110000000111110    1110000000111111    1110000001000000    1110000001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57405 - 57409

  --1110000001000010    1110000001000011    1110000001000100    1110000001000101    1110000001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57410 - 57414

  --1110000001000111    1110000001001000    1110000001001001    1110000001001010    1110000001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57415 - 57419

  --1110000001001100    1110000001001101    1110000001001110    1110000001001111    1110000001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57420 - 57424

  --1110000001010001    1110000001010010    1110000001010011    1110000001010100    1110000001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57425 - 57429

  --1110000001010110    1110000001010111    1110000001011000    1110000001011001    1110000001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57430 - 57434

  --1110000001011011    1110000001011100    1110000001011101    1110000001011110    1110000001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57435 - 57439

  --1110000001100000    1110000001100001    1110000001100010    1110000001100011    1110000001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57440 - 57444

  --1110000001100101    1110000001100110    1110000001100111    1110000001101000    1110000001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57445 - 57449

  --1110000001101010    1110000001101011    1110000001101100    1110000001101101    1110000001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57450 - 57454

  --1110000001101111    1110000001110000    1110000001110001    1110000001110010    1110000001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57455 - 57459

  --1110000001110100    1110000001110101    1110000001110110    1110000001110111    1110000001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57460 - 57464

  --1110000001111001    1110000001111010    1110000001111011    1110000001111100    1110000001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57465 - 57469

  --1110000001111110    1110000001111111    1110000010000000    1110000010000001    1110000010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57470 - 57474

  --1110000010000011    1110000010000100    1110000010000101    1110000010000110    1110000010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57475 - 57479

  --1110000010001000    1110000010001001    1110000010001010    1110000010001011    1110000010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57480 - 57484

  --1110000010001101    1110000010001110    1110000010001111    1110000010010000    1110000010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57485 - 57489

  --1110000010010010    1110000010010011    1110000010010100    1110000010010101    1110000010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57490 - 57494

  --1110000010010111    1110000010011000    1110000010011001    1110000010011010    1110000010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57495 - 57499

  --1110000010011100    1110000010011101    1110000010011110    1110000010011111    1110000010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57500 - 57504

  --1110000010100001    1110000010100010    1110000010100011    1110000010100100    1110000010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57505 - 57509

  --1110000010100110    1110000010100111    1110000010101000    1110000010101001    1110000010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57510 - 57514

  --1110000010101011    1110000010101100    1110000010101101    1110000010101110    1110000010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57515 - 57519

  --1110000010110000    1110000010110001    1110000010110010    1110000010110011    1110000010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57520 - 57524

  --1110000010110101    1110000010110110    1110000010110111    1110000010111000    1110000010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57525 - 57529

  --1110000010111010    1110000010111011    1110000010111100    1110000010111101    1110000010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57530 - 57534

  --1110000010111111    1110000011000000    1110000011000001    1110000011000010    1110000011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57535 - 57539

  --1110000011000100    1110000011000101    1110000011000110    1110000011000111    1110000011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57540 - 57544

  --1110000011001001    1110000011001010    1110000011001011    1110000011001100    1110000011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57545 - 57549

  --1110000011001110    1110000011001111    1110000011010000    1110000011010001    1110000011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57550 - 57554

  --1110000011010011    1110000011010100    1110000011010101    1110000011010110    1110000011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57555 - 57559

  --1110000011011000    1110000011011001    1110000011011010    1110000011011011    1110000011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57560 - 57564

  --1110000011011101    1110000011011110    1110000011011111    1110000011100000    1110000011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57565 - 57569

  --1110000011100010    1110000011100011    1110000011100100    1110000011100101    1110000011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57570 - 57574

  --1110000011100111    1110000011101000    1110000011101001    1110000011101010    1110000011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57575 - 57579

  --1110000011101100    1110000011101101    1110000011101110    1110000011101111    1110000011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57580 - 57584

  --1110000011110001    1110000011110010    1110000011110011    1110000011110100    1110000011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57585 - 57589

  --1110000011110110    1110000011110111    1110000011111000    1110000011111001    1110000011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57590 - 57594

  --1110000011111011    1110000011111100    1110000011111101    1110000011111110    1110000011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57595 - 57599

  --1110000100000000    1110000100000001    1110000100000010    1110000100000011    1110000100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57600 - 57604

  --1110000100000101    1110000100000110    1110000100000111    1110000100001000    1110000100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57605 - 57609

  --1110000100001010    1110000100001011    1110000100001100    1110000100001101    1110000100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57610 - 57614

  --1110000100001111    1110000100010000    1110000100010001    1110000100010010    1110000100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57615 - 57619

  --1110000100010100    1110000100010101    1110000100010110    1110000100010111    1110000100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57620 - 57624

  --1110000100011001    1110000100011010    1110000100011011    1110000100011100    1110000100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57625 - 57629

  --1110000100011110    1110000100011111    1110000100100000    1110000100100001    1110000100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57630 - 57634

  --1110000100100011    1110000100100100    1110000100100101    1110000100100110    1110000100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57635 - 57639

  --1110000100101000    1110000100101001    1110000100101010    1110000100101011    1110000100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57640 - 57644

  --1110000100101101    1110000100101110    1110000100101111    1110000100110000    1110000100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57645 - 57649

  --1110000100110010    1110000100110011    1110000100110100    1110000100110101    1110000100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57650 - 57654

  --1110000100110111    1110000100111000    1110000100111001    1110000100111010    1110000100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57655 - 57659

  --1110000100111100    1110000100111101    1110000100111110    1110000100111111    1110000101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57660 - 57664

  --1110000101000001    1110000101000010    1110000101000011    1110000101000100    1110000101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57665 - 57669

  --1110000101000110    1110000101000111    1110000101001000    1110000101001001    1110000101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57670 - 57674

  --1110000101001011    1110000101001100    1110000101001101    1110000101001110    1110000101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57675 - 57679

  --1110000101010000    1110000101010001    1110000101010010    1110000101010011    1110000101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57680 - 57684

  --1110000101010101    1110000101010110    1110000101010111    1110000101011000    1110000101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57685 - 57689

  --1110000101011010    1110000101011011    1110000101011100    1110000101011101    1110000101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57690 - 57694

  --1110000101011111    1110000101100000    1110000101100001    1110000101100010    1110000101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57695 - 57699

  --1110000101100100    1110000101100101    1110000101100110    1110000101100111    1110000101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57700 - 57704

  --1110000101101001    1110000101101010    1110000101101011    1110000101101100    1110000101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57705 - 57709

  --1110000101101110    1110000101101111    1110000101110000    1110000101110001    1110000101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57710 - 57714

  --1110000101110011    1110000101110100    1110000101110101    1110000101110110    1110000101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57715 - 57719

  --1110000101111000    1110000101111001    1110000101111010    1110000101111011    1110000101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57720 - 57724

  --1110000101111101    1110000101111110    1110000101111111    1110000110000000    1110000110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57725 - 57729

  --1110000110000010    1110000110000011    1110000110000100    1110000110000101    1110000110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57730 - 57734

  --1110000110000111    1110000110001000    1110000110001001    1110000110001010    1110000110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57735 - 57739

  --1110000110001100    1110000110001101    1110000110001110    1110000110001111    1110000110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57740 - 57744

  --1110000110010001    1110000110010010    1110000110010011    1110000110010100    1110000110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57745 - 57749

  --1110000110010110    1110000110010111    1110000110011000    1110000110011001    1110000110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57750 - 57754

  --1110000110011011    1110000110011100    1110000110011101    1110000110011110    1110000110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57755 - 57759

  --1110000110100000    1110000110100001    1110000110100010    1110000110100011    1110000110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57760 - 57764

  --1110000110100101    1110000110100110    1110000110100111    1110000110101000    1110000110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57765 - 57769

  --1110000110101010    1110000110101011    1110000110101100    1110000110101101    1110000110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57770 - 57774

  --1110000110101111    1110000110110000    1110000110110001    1110000110110010    1110000110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57775 - 57779

  --1110000110110100    1110000110110101    1110000110110110    1110000110110111    1110000110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57780 - 57784

  --1110000110111001    1110000110111010    1110000110111011    1110000110111100    1110000110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57785 - 57789

  --1110000110111110    1110000110111111    1110000111000000    1110000111000001    1110000111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57790 - 57794

  --1110000111000011    1110000111000100    1110000111000101    1110000111000110    1110000111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57795 - 57799

  --1110000111001000    1110000111001001    1110000111001010    1110000111001011    1110000111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57800 - 57804

  --1110000111001101    1110000111001110    1110000111001111    1110000111010000    1110000111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57805 - 57809

  --1110000111010010    1110000111010011    1110000111010100    1110000111010101    1110000111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57810 - 57814

  --1110000111010111    1110000111011000    1110000111011001    1110000111011010    1110000111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57815 - 57819

  --1110000111011100    1110000111011101    1110000111011110    1110000111011111    1110000111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57820 - 57824

  --1110000111100001    1110000111100010    1110000111100011    1110000111100100    1110000111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57825 - 57829

  --1110000111100110    1110000111100111    1110000111101000    1110000111101001    1110000111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57830 - 57834

  --1110000111101011    1110000111101100    1110000111101101    1110000111101110    1110000111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57835 - 57839

  --1110000111110000    1110000111110001    1110000111110010    1110000111110011    1110000111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57840 - 57844

  --1110000111110101    1110000111110110    1110000111110111    1110000111111000    1110000111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57845 - 57849

  --1110000111111010    1110000111111011    1110000111111100    1110000111111101    1110000111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57850 - 57854

  --1110000111111111    1110001000000000    1110001000000001    1110001000000010    1110001000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57855 - 57859

  --1110001000000100    1110001000000101    1110001000000110    1110001000000111    1110001000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57860 - 57864

  --1110001000001001    1110001000001010    1110001000001011    1110001000001100    1110001000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57865 - 57869

  --1110001000001110    1110001000001111    1110001000010000    1110001000010001    1110001000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57870 - 57874

  --1110001000010011    1110001000010100    1110001000010101    1110001000010110    1110001000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57875 - 57879

  --1110001000011000    1110001000011001    1110001000011010    1110001000011011    1110001000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57880 - 57884

  --1110001000011101    1110001000011110    1110001000011111    1110001000100000    1110001000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57885 - 57889

  --1110001000100010    1110001000100011    1110001000100100    1110001000100101    1110001000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57890 - 57894

  --1110001000100111    1110001000101000    1110001000101001    1110001000101010    1110001000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57895 - 57899

  --1110001000101100    1110001000101101    1110001000101110    1110001000101111    1110001000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57900 - 57904

  --1110001000110001    1110001000110010    1110001000110011    1110001000110100    1110001000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57905 - 57909

  --1110001000110110    1110001000110111    1110001000111000    1110001000111001    1110001000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57910 - 57914

  --1110001000111011    1110001000111100    1110001000111101    1110001000111110    1110001000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57915 - 57919

  --1110001001000000    1110001001000001    1110001001000010    1110001001000011    1110001001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57920 - 57924

  --1110001001000101    1110001001000110    1110001001000111    1110001001001000    1110001001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57925 - 57929

  --1110001001001010    1110001001001011    1110001001001100    1110001001001101    1110001001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57930 - 57934

  --1110001001001111    1110001001010000    1110001001010001    1110001001010010    1110001001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57935 - 57939

  --1110001001010100    1110001001010101    1110001001010110    1110001001010111    1110001001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57940 - 57944

  --1110001001011001    1110001001011010    1110001001011011    1110001001011100    1110001001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57945 - 57949

  --1110001001011110    1110001001011111    1110001001100000    1110001001100001    1110001001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57950 - 57954

  --1110001001100011    1110001001100100    1110001001100101    1110001001100110    1110001001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57955 - 57959

  --1110001001101000    1110001001101001    1110001001101010    1110001001101011    1110001001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57960 - 57964

  --1110001001101101    1110001001101110    1110001001101111    1110001001110000    1110001001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57965 - 57969

  --1110001001110010    1110001001110011    1110001001110100    1110001001110101    1110001001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57970 - 57974

  --1110001001110111    1110001001111000    1110001001111001    1110001001111010    1110001001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57975 - 57979

  --1110001001111100    1110001001111101    1110001001111110    1110001001111111    1110001010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57980 - 57984

  --1110001010000001    1110001010000010    1110001010000011    1110001010000100    1110001010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57985 - 57989

  --1110001010000110    1110001010000111    1110001010001000    1110001010001001    1110001010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57990 - 57994

  --1110001010001011    1110001010001100    1110001010001101    1110001010001110    1110001010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 57995 - 57999

  --1110001010010000    1110001010010001    1110001010010010    1110001010010011    1110001010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58000 - 58004

  --1110001010010101    1110001010010110    1110001010010111    1110001010011000    1110001010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58005 - 58009

  --1110001010011010    1110001010011011    1110001010011100    1110001010011101    1110001010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58010 - 58014

  --1110001010011111    1110001010100000    1110001010100001    1110001010100010    1110001010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58015 - 58019

  --1110001010100100    1110001010100101    1110001010100110    1110001010100111    1110001010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58020 - 58024

  --1110001010101001    1110001010101010    1110001010101011    1110001010101100    1110001010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58025 - 58029

  --1110001010101110    1110001010101111    1110001010110000    1110001010110001    1110001010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58030 - 58034

  --1110001010110011    1110001010110100    1110001010110101    1110001010110110    1110001010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58035 - 58039

  --1110001010111000    1110001010111001    1110001010111010    1110001010111011    1110001010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58040 - 58044

  --1110001010111101    1110001010111110    1110001010111111    1110001011000000    1110001011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58045 - 58049

  --1110001011000010    1110001011000011    1110001011000100    1110001011000101    1110001011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58050 - 58054

  --1110001011000111    1110001011001000    1110001011001001    1110001011001010    1110001011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58055 - 58059

  --1110001011001100    1110001011001101    1110001011001110    1110001011001111    1110001011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58060 - 58064

  --1110001011010001    1110001011010010    1110001011010011    1110001011010100    1110001011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58065 - 58069

  --1110001011010110    1110001011010111    1110001011011000    1110001011011001    1110001011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58070 - 58074

  --1110001011011011    1110001011011100    1110001011011101    1110001011011110    1110001011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58075 - 58079

  --1110001011100000    1110001011100001    1110001011100010    1110001011100011    1110001011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58080 - 58084

  --1110001011100101    1110001011100110    1110001011100111    1110001011101000    1110001011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58085 - 58089

  --1110001011101010    1110001011101011    1110001011101100    1110001011101101    1110001011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58090 - 58094

  --1110001011101111    1110001011110000    1110001011110001    1110001011110010    1110001011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58095 - 58099

  --1110001011110100    1110001011110101    1110001011110110    1110001011110111    1110001011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58100 - 58104

  --1110001011111001    1110001011111010    1110001011111011    1110001011111100    1110001011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58105 - 58109

  --1110001011111110    1110001011111111    1110001100000000    1110001100000001    1110001100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58110 - 58114

  --1110001100000011    1110001100000100    1110001100000101    1110001100000110    1110001100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58115 - 58119

  --1110001100001000    1110001100001001    1110001100001010    1110001100001011    1110001100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58120 - 58124

  --1110001100001101    1110001100001110    1110001100001111    1110001100010000    1110001100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58125 - 58129

  --1110001100010010    1110001100010011    1110001100010100    1110001100010101    1110001100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58130 - 58134

  --1110001100010111    1110001100011000    1110001100011001    1110001100011010    1110001100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58135 - 58139

  --1110001100011100    1110001100011101    1110001100011110    1110001100011111    1110001100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58140 - 58144

  --1110001100100001    1110001100100010    1110001100100011    1110001100100100    1110001100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58145 - 58149

  --1110001100100110    1110001100100111    1110001100101000    1110001100101001    1110001100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58150 - 58154

  --1110001100101011    1110001100101100    1110001100101101    1110001100101110    1110001100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58155 - 58159

  --1110001100110000    1110001100110001    1110001100110010    1110001100110011    1110001100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58160 - 58164

  --1110001100110101    1110001100110110    1110001100110111    1110001100111000    1110001100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58165 - 58169

  --1110001100111010    1110001100111011    1110001100111100    1110001100111101    1110001100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58170 - 58174

  --1110001100111111    1110001101000000    1110001101000001    1110001101000010    1110001101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58175 - 58179

  --1110001101000100    1110001101000101    1110001101000110    1110001101000111    1110001101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58180 - 58184

  --1110001101001001    1110001101001010    1110001101001011    1110001101001100    1110001101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58185 - 58189

  --1110001101001110    1110001101001111    1110001101010000    1110001101010001    1110001101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58190 - 58194

  --1110001101010011    1110001101010100    1110001101010101    1110001101010110    1110001101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58195 - 58199

  --1110001101011000    1110001101011001    1110001101011010    1110001101011011    1110001101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58200 - 58204

  --1110001101011101    1110001101011110    1110001101011111    1110001101100000    1110001101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58205 - 58209

  --1110001101100010    1110001101100011    1110001101100100    1110001101100101    1110001101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58210 - 58214

  --1110001101100111    1110001101101000    1110001101101001    1110001101101010    1110001101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58215 - 58219

  --1110001101101100    1110001101101101    1110001101101110    1110001101101111    1110001101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58220 - 58224

  --1110001101110001    1110001101110010    1110001101110011    1110001101110100    1110001101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58225 - 58229

  --1110001101110110    1110001101110111    1110001101111000    1110001101111001    1110001101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58230 - 58234

  --1110001101111011    1110001101111100    1110001101111101    1110001101111110    1110001101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58235 - 58239

  --1110001110000000    1110001110000001    1110001110000010    1110001110000011    1110001110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58240 - 58244

  --1110001110000101    1110001110000110    1110001110000111    1110001110001000    1110001110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58245 - 58249

  --1110001110001010    1110001110001011    1110001110001100    1110001110001101    1110001110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58250 - 58254

  --1110001110001111    1110001110010000    1110001110010001    1110001110010010    1110001110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58255 - 58259

  --1110001110010100    1110001110010101    1110001110010110    1110001110010111    1110001110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58260 - 58264

  --1110001110011001    1110001110011010    1110001110011011    1110001110011100    1110001110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58265 - 58269

  --1110001110011110    1110001110011111    1110001110100000    1110001110100001    1110001110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58270 - 58274

  --1110001110100011    1110001110100100    1110001110100101    1110001110100110    1110001110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58275 - 58279

  --1110001110101000    1110001110101001    1110001110101010    1110001110101011    1110001110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58280 - 58284

  --1110001110101101    1110001110101110    1110001110101111    1110001110110000    1110001110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58285 - 58289

  --1110001110110010    1110001110110011    1110001110110100    1110001110110101    1110001110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58290 - 58294

  --1110001110110111    1110001110111000    1110001110111001    1110001110111010    1110001110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58295 - 58299

  --1110001110111100    1110001110111101    1110001110111110    1110001110111111    1110001111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58300 - 58304

  --1110001111000001    1110001111000010    1110001111000011    1110001111000100    1110001111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58305 - 58309

  --1110001111000110    1110001111000111    1110001111001000    1110001111001001    1110001111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58310 - 58314

  --1110001111001011    1110001111001100    1110001111001101    1110001111001110    1110001111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58315 - 58319

  --1110001111010000    1110001111010001    1110001111010010    1110001111010011    1110001111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58320 - 58324

  --1110001111010101    1110001111010110    1110001111010111    1110001111011000    1110001111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58325 - 58329

  --1110001111011010    1110001111011011    1110001111011100    1110001111011101    1110001111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58330 - 58334

  --1110001111011111    1110001111100000    1110001111100001    1110001111100010    1110001111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58335 - 58339

  --1110001111100100    1110001111100101    1110001111100110    1110001111100111    1110001111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58340 - 58344

  --1110001111101001    1110001111101010    1110001111101011    1110001111101100    1110001111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58345 - 58349

  --1110001111101110    1110001111101111    1110001111110000    1110001111110001    1110001111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58350 - 58354

  --1110001111110011    1110001111110100    1110001111110101    1110001111110110    1110001111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58355 - 58359

  --1110001111111000    1110001111111001    1110001111111010    1110001111111011    1110001111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58360 - 58364

  --1110001111111101    1110001111111110    1110001111111111    1110010000000000    1110010000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58365 - 58369

  --1110010000000010    1110010000000011    1110010000000100    1110010000000101    1110010000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58370 - 58374

  --1110010000000111    1110010000001000    1110010000001001    1110010000001010    1110010000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58375 - 58379

  --1110010000001100    1110010000001101    1110010000001110    1110010000001111    1110010000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58380 - 58384

  --1110010000010001    1110010000010010    1110010000010011    1110010000010100    1110010000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58385 - 58389

  --1110010000010110    1110010000010111    1110010000011000    1110010000011001    1110010000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58390 - 58394

  --1110010000011011    1110010000011100    1110010000011101    1110010000011110    1110010000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58395 - 58399

  --1110010000100000    1110010000100001    1110010000100010    1110010000100011    1110010000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58400 - 58404

  --1110010000100101    1110010000100110    1110010000100111    1110010000101000    1110010000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58405 - 58409

  --1110010000101010    1110010000101011    1110010000101100    1110010000101101    1110010000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58410 - 58414

  --1110010000101111    1110010000110000    1110010000110001    1110010000110010    1110010000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58415 - 58419

  --1110010000110100    1110010000110101    1110010000110110    1110010000110111    1110010000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58420 - 58424

  --1110010000111001    1110010000111010    1110010000111011    1110010000111100    1110010000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58425 - 58429

  --1110010000111110    1110010000111111    1110010001000000    1110010001000001    1110010001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58430 - 58434

  --1110010001000011    1110010001000100    1110010001000101    1110010001000110    1110010001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58435 - 58439

  --1110010001001000    1110010001001001    1110010001001010    1110010001001011    1110010001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58440 - 58444

  --1110010001001101    1110010001001110    1110010001001111    1110010001010000    1110010001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58445 - 58449

  --1110010001010010    1110010001010011    1110010001010100    1110010001010101    1110010001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58450 - 58454

  --1110010001010111    1110010001011000    1110010001011001    1110010001011010    1110010001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58455 - 58459

  --1110010001011100    1110010001011101    1110010001011110    1110010001011111    1110010001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58460 - 58464

  --1110010001100001    1110010001100010    1110010001100011    1110010001100100    1110010001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58465 - 58469

  --1110010001100110    1110010001100111    1110010001101000    1110010001101001    1110010001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58470 - 58474

  --1110010001101011    1110010001101100    1110010001101101    1110010001101110    1110010001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58475 - 58479

  --1110010001110000    1110010001110001    1110010001110010    1110010001110011    1110010001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58480 - 58484

  --1110010001110101    1110010001110110    1110010001110111    1110010001111000    1110010001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58485 - 58489

  --1110010001111010    1110010001111011    1110010001111100    1110010001111101    1110010001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58490 - 58494

  --1110010001111111    1110010010000000    1110010010000001    1110010010000010    1110010010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58495 - 58499

  --1110010010000100    1110010010000101    1110010010000110    1110010010000111    1110010010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58500 - 58504

  --1110010010001001    1110010010001010    1110010010001011    1110010010001100    1110010010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58505 - 58509

  --1110010010001110    1110010010001111    1110010010010000    1110010010010001    1110010010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58510 - 58514

  --1110010010010011    1110010010010100    1110010010010101    1110010010010110    1110010010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58515 - 58519

  --1110010010011000    1110010010011001    1110010010011010    1110010010011011    1110010010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58520 - 58524

  --1110010010011101    1110010010011110    1110010010011111    1110010010100000    1110010010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58525 - 58529

  --1110010010100010    1110010010100011    1110010010100100    1110010010100101    1110010010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58530 - 58534

  --1110010010100111    1110010010101000    1110010010101001    1110010010101010    1110010010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58535 - 58539

  --1110010010101100    1110010010101101    1110010010101110    1110010010101111    1110010010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58540 - 58544

  --1110010010110001    1110010010110010    1110010010110011    1110010010110100    1110010010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58545 - 58549

  --1110010010110110    1110010010110111    1110010010111000    1110010010111001    1110010010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58550 - 58554

  --1110010010111011    1110010010111100    1110010010111101    1110010010111110    1110010010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58555 - 58559

  --1110010011000000    1110010011000001    1110010011000010    1110010011000011    1110010011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58560 - 58564

  --1110010011000101    1110010011000110    1110010011000111    1110010011001000    1110010011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58565 - 58569

  --1110010011001010    1110010011001011    1110010011001100    1110010011001101    1110010011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58570 - 58574

  --1110010011001111    1110010011010000    1110010011010001    1110010011010010    1110010011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58575 - 58579

  --1110010011010100    1110010011010101    1110010011010110    1110010011010111    1110010011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58580 - 58584

  --1110010011011001    1110010011011010    1110010011011011    1110010011011100    1110010011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58585 - 58589

  --1110010011011110    1110010011011111    1110010011100000    1110010011100001    1110010011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58590 - 58594

  --1110010011100011    1110010011100100    1110010011100101    1110010011100110    1110010011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58595 - 58599

  --1110010011101000    1110010011101001    1110010011101010    1110010011101011    1110010011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58600 - 58604

  --1110010011101101    1110010011101110    1110010011101111    1110010011110000    1110010011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58605 - 58609

  --1110010011110010    1110010011110011    1110010011110100    1110010011110101    1110010011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58610 - 58614

  --1110010011110111    1110010011111000    1110010011111001    1110010011111010    1110010011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58615 - 58619

  --1110010011111100    1110010011111101    1110010011111110    1110010011111111    1110010100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58620 - 58624

  --1110010100000001    1110010100000010    1110010100000011    1110010100000100    1110010100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58625 - 58629

  --1110010100000110    1110010100000111    1110010100001000    1110010100001001    1110010100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58630 - 58634

  --1110010100001011    1110010100001100    1110010100001101    1110010100001110    1110010100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58635 - 58639

  --1110010100010000    1110010100010001    1110010100010010    1110010100010011    1110010100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58640 - 58644

  --1110010100010101    1110010100010110    1110010100010111    1110010100011000    1110010100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58645 - 58649

  --1110010100011010    1110010100011011    1110010100011100    1110010100011101    1110010100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58650 - 58654

  --1110010100011111    1110010100100000    1110010100100001    1110010100100010    1110010100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58655 - 58659

  --1110010100100100    1110010100100101    1110010100100110    1110010100100111    1110010100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58660 - 58664

  --1110010100101001    1110010100101010    1110010100101011    1110010100101100    1110010100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58665 - 58669

  --1110010100101110    1110010100101111    1110010100110000    1110010100110001    1110010100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58670 - 58674

  --1110010100110011    1110010100110100    1110010100110101    1110010100110110    1110010100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58675 - 58679

  --1110010100111000    1110010100111001    1110010100111010    1110010100111011    1110010100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58680 - 58684

  --1110010100111101    1110010100111110    1110010100111111    1110010101000000    1110010101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58685 - 58689

  --1110010101000010    1110010101000011    1110010101000100    1110010101000101    1110010101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58690 - 58694

  --1110010101000111    1110010101001000    1110010101001001    1110010101001010    1110010101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58695 - 58699

  --1110010101001100    1110010101001101    1110010101001110    1110010101001111    1110010101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58700 - 58704

  --1110010101010001    1110010101010010    1110010101010011    1110010101010100    1110010101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58705 - 58709

  --1110010101010110    1110010101010111    1110010101011000    1110010101011001    1110010101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58710 - 58714

  --1110010101011011    1110010101011100    1110010101011101    1110010101011110    1110010101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58715 - 58719

  --1110010101100000    1110010101100001    1110010101100010    1110010101100011    1110010101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58720 - 58724

  --1110010101100101    1110010101100110    1110010101100111    1110010101101000    1110010101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58725 - 58729

  --1110010101101010    1110010101101011    1110010101101100    1110010101101101    1110010101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58730 - 58734

  --1110010101101111    1110010101110000    1110010101110001    1110010101110010    1110010101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58735 - 58739

  --1110010101110100    1110010101110101    1110010101110110    1110010101110111    1110010101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58740 - 58744

  --1110010101111001    1110010101111010    1110010101111011    1110010101111100    1110010101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58745 - 58749

  --1110010101111110    1110010101111111    1110010110000000    1110010110000001    1110010110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58750 - 58754

  --1110010110000011    1110010110000100    1110010110000101    1110010110000110    1110010110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58755 - 58759

  --1110010110001000    1110010110001001    1110010110001010    1110010110001011    1110010110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58760 - 58764

  --1110010110001101    1110010110001110    1110010110001111    1110010110010000    1110010110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58765 - 58769

  --1110010110010010    1110010110010011    1110010110010100    1110010110010101    1110010110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58770 - 58774

  --1110010110010111    1110010110011000    1110010110011001    1110010110011010    1110010110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58775 - 58779

  --1110010110011100    1110010110011101    1110010110011110    1110010110011111    1110010110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58780 - 58784

  --1110010110100001    1110010110100010    1110010110100011    1110010110100100    1110010110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58785 - 58789

  --1110010110100110    1110010110100111    1110010110101000    1110010110101001    1110010110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58790 - 58794

  --1110010110101011    1110010110101100    1110010110101101    1110010110101110    1110010110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58795 - 58799

  --1110010110110000    1110010110110001    1110010110110010    1110010110110011    1110010110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58800 - 58804

  --1110010110110101    1110010110110110    1110010110110111    1110010110111000    1110010110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58805 - 58809

  --1110010110111010    1110010110111011    1110010110111100    1110010110111101    1110010110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58810 - 58814

  --1110010110111111    1110010111000000    1110010111000001    1110010111000010    1110010111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58815 - 58819

  --1110010111000100    1110010111000101    1110010111000110    1110010111000111    1110010111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58820 - 58824

  --1110010111001001    1110010111001010    1110010111001011    1110010111001100    1110010111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58825 - 58829

  --1110010111001110    1110010111001111    1110010111010000    1110010111010001    1110010111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58830 - 58834

  --1110010111010011    1110010111010100    1110010111010101    1110010111010110    1110010111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58835 - 58839

  --1110010111011000    1110010111011001    1110010111011010    1110010111011011    1110010111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58840 - 58844

  --1110010111011101    1110010111011110    1110010111011111    1110010111100000    1110010111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58845 - 58849

  --1110010111100010    1110010111100011    1110010111100100    1110010111100101    1110010111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58850 - 58854

  --1110010111100111    1110010111101000    1110010111101001    1110010111101010    1110010111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58855 - 58859

  --1110010111101100    1110010111101101    1110010111101110    1110010111101111    1110010111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58860 - 58864

  --1110010111110001    1110010111110010    1110010111110011    1110010111110100    1110010111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58865 - 58869

  --1110010111110110    1110010111110111    1110010111111000    1110010111111001    1110010111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58870 - 58874

  --1110010111111011    1110010111111100    1110010111111101    1110010111111110    1110010111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58875 - 58879

  --1110011000000000    1110011000000001    1110011000000010    1110011000000011    1110011000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58880 - 58884

  --1110011000000101    1110011000000110    1110011000000111    1110011000001000    1110011000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58885 - 58889

  --1110011000001010    1110011000001011    1110011000001100    1110011000001101    1110011000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58890 - 58894

  --1110011000001111    1110011000010000    1110011000010001    1110011000010010    1110011000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58895 - 58899

  --1110011000010100    1110011000010101    1110011000010110    1110011000010111    1110011000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58900 - 58904

  --1110011000011001    1110011000011010    1110011000011011    1110011000011100    1110011000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58905 - 58909

  --1110011000011110    1110011000011111    1110011000100000    1110011000100001    1110011000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58910 - 58914

  --1110011000100011    1110011000100100    1110011000100101    1110011000100110    1110011000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58915 - 58919

  --1110011000101000    1110011000101001    1110011000101010    1110011000101011    1110011000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58920 - 58924

  --1110011000101101    1110011000101110    1110011000101111    1110011000110000    1110011000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58925 - 58929

  --1110011000110010    1110011000110011    1110011000110100    1110011000110101    1110011000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58930 - 58934

  --1110011000110111    1110011000111000    1110011000111001    1110011000111010    1110011000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58935 - 58939

  --1110011000111100    1110011000111101    1110011000111110    1110011000111111    1110011001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58940 - 58944

  --1110011001000001    1110011001000010    1110011001000011    1110011001000100    1110011001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58945 - 58949

  --1110011001000110    1110011001000111    1110011001001000    1110011001001001    1110011001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58950 - 58954

  --1110011001001011    1110011001001100    1110011001001101    1110011001001110    1110011001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58955 - 58959

  --1110011001010000    1110011001010001    1110011001010010    1110011001010011    1110011001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58960 - 58964

  --1110011001010101    1110011001010110    1110011001010111    1110011001011000    1110011001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58965 - 58969

  --1110011001011010    1110011001011011    1110011001011100    1110011001011101    1110011001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58970 - 58974

  --1110011001011111    1110011001100000    1110011001100001    1110011001100010    1110011001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58975 - 58979

  --1110011001100100    1110011001100101    1110011001100110    1110011001100111    1110011001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58980 - 58984

  --1110011001101001    1110011001101010    1110011001101011    1110011001101100    1110011001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58985 - 58989

  --1110011001101110    1110011001101111    1110011001110000    1110011001110001    1110011001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58990 - 58994

  --1110011001110011    1110011001110100    1110011001110101    1110011001110110    1110011001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 58995 - 58999

  --1110011001111000    1110011001111001    1110011001111010    1110011001111011    1110011001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59000 - 59004

  --1110011001111101    1110011001111110    1110011001111111    1110011010000000    1110011010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59005 - 59009

  --1110011010000010    1110011010000011    1110011010000100    1110011010000101    1110011010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59010 - 59014

  --1110011010000111    1110011010001000    1110011010001001    1110011010001010    1110011010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59015 - 59019

  --1110011010001100    1110011010001101    1110011010001110    1110011010001111    1110011010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59020 - 59024

  --1110011010010001    1110011010010010    1110011010010011    1110011010010100    1110011010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59025 - 59029

  --1110011010010110    1110011010010111    1110011010011000    1110011010011001    1110011010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59030 - 59034

  --1110011010011011    1110011010011100    1110011010011101    1110011010011110    1110011010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59035 - 59039

  --1110011010100000    1110011010100001    1110011010100010    1110011010100011    1110011010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59040 - 59044

  --1110011010100101    1110011010100110    1110011010100111    1110011010101000    1110011010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59045 - 59049

  --1110011010101010    1110011010101011    1110011010101100    1110011010101101    1110011010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59050 - 59054

  --1110011010101111    1110011010110000    1110011010110001    1110011010110010    1110011010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59055 - 59059

  --1110011010110100    1110011010110101    1110011010110110    1110011010110111    1110011010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59060 - 59064

  --1110011010111001    1110011010111010    1110011010111011    1110011010111100    1110011010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59065 - 59069

  --1110011010111110    1110011010111111    1110011011000000    1110011011000001    1110011011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59070 - 59074

  --1110011011000011    1110011011000100    1110011011000101    1110011011000110    1110011011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59075 - 59079

  --1110011011001000    1110011011001001    1110011011001010    1110011011001011    1110011011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59080 - 59084

  --1110011011001101    1110011011001110    1110011011001111    1110011011010000    1110011011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59085 - 59089

  --1110011011010010    1110011011010011    1110011011010100    1110011011010101    1110011011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59090 - 59094

  --1110011011010111    1110011011011000    1110011011011001    1110011011011010    1110011011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59095 - 59099

  --1110011011011100    1110011011011101    1110011011011110    1110011011011111    1110011011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59100 - 59104

  --1110011011100001    1110011011100010    1110011011100011    1110011011100100    1110011011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59105 - 59109

  --1110011011100110    1110011011100111    1110011011101000    1110011011101001    1110011011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59110 - 59114

  --1110011011101011    1110011011101100    1110011011101101    1110011011101110    1110011011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59115 - 59119

  --1110011011110000    1110011011110001    1110011011110010    1110011011110011    1110011011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59120 - 59124

  --1110011011110101    1110011011110110    1110011011110111    1110011011111000    1110011011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59125 - 59129

  --1110011011111010    1110011011111011    1110011011111100    1110011011111101    1110011011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59130 - 59134

  --1110011011111111    1110011100000000    1110011100000001    1110011100000010    1110011100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59135 - 59139

  --1110011100000100    1110011100000101    1110011100000110    1110011100000111    1110011100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59140 - 59144

  --1110011100001001    1110011100001010    1110011100001011    1110011100001100    1110011100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59145 - 59149

  --1110011100001110    1110011100001111    1110011100010000    1110011100010001    1110011100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59150 - 59154

  --1110011100010011    1110011100010100    1110011100010101    1110011100010110    1110011100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59155 - 59159

  --1110011100011000    1110011100011001    1110011100011010    1110011100011011    1110011100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59160 - 59164

  --1110011100011101    1110011100011110    1110011100011111    1110011100100000    1110011100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59165 - 59169

  --1110011100100010    1110011100100011    1110011100100100    1110011100100101    1110011100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59170 - 59174

  --1110011100100111    1110011100101000    1110011100101001    1110011100101010    1110011100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59175 - 59179

  --1110011100101100    1110011100101101    1110011100101110    1110011100101111    1110011100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59180 - 59184

  --1110011100110001    1110011100110010    1110011100110011    1110011100110100    1110011100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59185 - 59189

  --1110011100110110    1110011100110111    1110011100111000    1110011100111001    1110011100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59190 - 59194

  --1110011100111011    1110011100111100    1110011100111101    1110011100111110    1110011100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59195 - 59199

  --1110011101000000    1110011101000001    1110011101000010    1110011101000011    1110011101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59200 - 59204

  --1110011101000101    1110011101000110    1110011101000111    1110011101001000    1110011101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59205 - 59209

  --1110011101001010    1110011101001011    1110011101001100    1110011101001101    1110011101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59210 - 59214

  --1110011101001111    1110011101010000    1110011101010001    1110011101010010    1110011101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59215 - 59219

  --1110011101010100    1110011101010101    1110011101010110    1110011101010111    1110011101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59220 - 59224

  --1110011101011001    1110011101011010    1110011101011011    1110011101011100    1110011101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59225 - 59229

  --1110011101011110    1110011101011111    1110011101100000    1110011101100001    1110011101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59230 - 59234

  --1110011101100011    1110011101100100    1110011101100101    1110011101100110    1110011101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59235 - 59239

  --1110011101101000    1110011101101001    1110011101101010    1110011101101011    1110011101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59240 - 59244

  --1110011101101101    1110011101101110    1110011101101111    1110011101110000    1110011101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59245 - 59249

  --1110011101110010    1110011101110011    1110011101110100    1110011101110101    1110011101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59250 - 59254

  --1110011101110111    1110011101111000    1110011101111001    1110011101111010    1110011101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59255 - 59259

  --1110011101111100    1110011101111101    1110011101111110    1110011101111111    1110011110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59260 - 59264

  --1110011110000001    1110011110000010    1110011110000011    1110011110000100    1110011110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59265 - 59269

  --1110011110000110    1110011110000111    1110011110001000    1110011110001001    1110011110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59270 - 59274

  --1110011110001011    1110011110001100    1110011110001101    1110011110001110    1110011110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59275 - 59279

  --1110011110010000    1110011110010001    1110011110010010    1110011110010011    1110011110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59280 - 59284

  --1110011110010101    1110011110010110    1110011110010111    1110011110011000    1110011110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59285 - 59289

  --1110011110011010    1110011110011011    1110011110011100    1110011110011101    1110011110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59290 - 59294

  --1110011110011111    1110011110100000    1110011110100001    1110011110100010    1110011110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59295 - 59299

  --1110011110100100    1110011110100101    1110011110100110    1110011110100111    1110011110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59300 - 59304

  --1110011110101001    1110011110101010    1110011110101011    1110011110101100    1110011110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59305 - 59309

  --1110011110101110    1110011110101111    1110011110110000    1110011110110001    1110011110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59310 - 59314

  --1110011110110011    1110011110110100    1110011110110101    1110011110110110    1110011110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59315 - 59319

  --1110011110111000    1110011110111001    1110011110111010    1110011110111011    1110011110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59320 - 59324

  --1110011110111101    1110011110111110    1110011110111111    1110011111000000    1110011111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59325 - 59329

  --1110011111000010    1110011111000011    1110011111000100    1110011111000101    1110011111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59330 - 59334

  --1110011111000111    1110011111001000    1110011111001001    1110011111001010    1110011111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59335 - 59339

  --1110011111001100    1110011111001101    1110011111001110    1110011111001111    1110011111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59340 - 59344

  --1110011111010001    1110011111010010    1110011111010011    1110011111010100    1110011111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59345 - 59349

  --1110011111010110    1110011111010111    1110011111011000    1110011111011001    1110011111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59350 - 59354

  --1110011111011011    1110011111011100    1110011111011101    1110011111011110    1110011111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59355 - 59359

  --1110011111100000    1110011111100001    1110011111100010    1110011111100011    1110011111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59360 - 59364

  --1110011111100101    1110011111100110    1110011111100111    1110011111101000    1110011111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59365 - 59369

  --1110011111101010    1110011111101011    1110011111101100    1110011111101101    1110011111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59370 - 59374

  --1110011111101111    1110011111110000    1110011111110001    1110011111110010    1110011111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59375 - 59379

  --1110011111110100    1110011111110101    1110011111110110    1110011111110111    1110011111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59380 - 59384

  --1110011111111001    1110011111111010    1110011111111011    1110011111111100    1110011111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59385 - 59389

  --1110011111111110    1110011111111111    1110100000000000    1110100000000001    1110100000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59390 - 59394

  --1110100000000011    1110100000000100    1110100000000101    1110100000000110    1110100000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59395 - 59399

  --1110100000001000    1110100000001001    1110100000001010    1110100000001011    1110100000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59400 - 59404

  --1110100000001101    1110100000001110    1110100000001111    1110100000010000    1110100000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59405 - 59409

  --1110100000010010    1110100000010011    1110100000010100    1110100000010101    1110100000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59410 - 59414

  --1110100000010111    1110100000011000    1110100000011001    1110100000011010    1110100000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59415 - 59419

  --1110100000011100    1110100000011101    1110100000011110    1110100000011111    1110100000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59420 - 59424

  --1110100000100001    1110100000100010    1110100000100011    1110100000100100    1110100000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59425 - 59429

  --1110100000100110    1110100000100111    1110100000101000    1110100000101001    1110100000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59430 - 59434

  --1110100000101011    1110100000101100    1110100000101101    1110100000101110    1110100000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59435 - 59439

  --1110100000110000    1110100000110001    1110100000110010    1110100000110011    1110100000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59440 - 59444

  --1110100000110101    1110100000110110    1110100000110111    1110100000111000    1110100000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59445 - 59449

  --1110100000111010    1110100000111011    1110100000111100    1110100000111101    1110100000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59450 - 59454

  --1110100000111111    1110100001000000    1110100001000001    1110100001000010    1110100001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59455 - 59459

  --1110100001000100    1110100001000101    1110100001000110    1110100001000111    1110100001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59460 - 59464

  --1110100001001001    1110100001001010    1110100001001011    1110100001001100    1110100001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59465 - 59469

  --1110100001001110    1110100001001111    1110100001010000    1110100001010001    1110100001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59470 - 59474

  --1110100001010011    1110100001010100    1110100001010101    1110100001010110    1110100001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59475 - 59479

  --1110100001011000    1110100001011001    1110100001011010    1110100001011011    1110100001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59480 - 59484

  --1110100001011101    1110100001011110    1110100001011111    1110100001100000    1110100001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59485 - 59489

  --1110100001100010    1110100001100011    1110100001100100    1110100001100101    1110100001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59490 - 59494

  --1110100001100111    1110100001101000    1110100001101001    1110100001101010    1110100001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59495 - 59499

  --1110100001101100    1110100001101101    1110100001101110    1110100001101111    1110100001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59500 - 59504

  --1110100001110001    1110100001110010    1110100001110011    1110100001110100    1110100001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59505 - 59509

  --1110100001110110    1110100001110111    1110100001111000    1110100001111001    1110100001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59510 - 59514

  --1110100001111011    1110100001111100    1110100001111101    1110100001111110    1110100001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59515 - 59519

  --1110100010000000    1110100010000001    1110100010000010    1110100010000011    1110100010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59520 - 59524

  --1110100010000101    1110100010000110    1110100010000111    1110100010001000    1110100010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59525 - 59529

  --1110100010001010    1110100010001011    1110100010001100    1110100010001101    1110100010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59530 - 59534

  --1110100010001111    1110100010010000    1110100010010001    1110100010010010    1110100010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59535 - 59539

  --1110100010010100    1110100010010101    1110100010010110    1110100010010111    1110100010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59540 - 59544

  --1110100010011001    1110100010011010    1110100010011011    1110100010011100    1110100010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59545 - 59549

  --1110100010011110    1110100010011111    1110100010100000    1110100010100001    1110100010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59550 - 59554

  --1110100010100011    1110100010100100    1110100010100101    1110100010100110    1110100010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59555 - 59559

  --1110100010101000    1110100010101001    1110100010101010    1110100010101011    1110100010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59560 - 59564

  --1110100010101101    1110100010101110    1110100010101111    1110100010110000    1110100010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59565 - 59569

  --1110100010110010    1110100010110011    1110100010110100    1110100010110101    1110100010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59570 - 59574

  --1110100010110111    1110100010111000    1110100010111001    1110100010111010    1110100010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59575 - 59579

  --1110100010111100    1110100010111101    1110100010111110    1110100010111111    1110100011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59580 - 59584

  --1110100011000001    1110100011000010    1110100011000011    1110100011000100    1110100011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59585 - 59589

  --1110100011000110    1110100011000111    1110100011001000    1110100011001001    1110100011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59590 - 59594

  --1110100011001011    1110100011001100    1110100011001101    1110100011001110    1110100011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59595 - 59599

  --1110100011010000    1110100011010001    1110100011010010    1110100011010011    1110100011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59600 - 59604

  --1110100011010101    1110100011010110    1110100011010111    1110100011011000    1110100011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59605 - 59609

  --1110100011011010    1110100011011011    1110100011011100    1110100011011101    1110100011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59610 - 59614

  --1110100011011111    1110100011100000    1110100011100001    1110100011100010    1110100011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59615 - 59619

  --1110100011100100    1110100011100101    1110100011100110    1110100011100111    1110100011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59620 - 59624

  --1110100011101001    1110100011101010    1110100011101011    1110100011101100    1110100011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59625 - 59629

  --1110100011101110    1110100011101111    1110100011110000    1110100011110001    1110100011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59630 - 59634

  --1110100011110011    1110100011110100    1110100011110101    1110100011110110    1110100011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59635 - 59639

  --1110100011111000    1110100011111001    1110100011111010    1110100011111011    1110100011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59640 - 59644

  --1110100011111101    1110100011111110    1110100011111111    1110100100000000    1110100100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59645 - 59649

  --1110100100000010    1110100100000011    1110100100000100    1110100100000101    1110100100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59650 - 59654

  --1110100100000111    1110100100001000    1110100100001001    1110100100001010    1110100100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59655 - 59659

  --1110100100001100    1110100100001101    1110100100001110    1110100100001111    1110100100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59660 - 59664

  --1110100100010001    1110100100010010    1110100100010011    1110100100010100    1110100100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59665 - 59669

  --1110100100010110    1110100100010111    1110100100011000    1110100100011001    1110100100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59670 - 59674

  --1110100100011011    1110100100011100    1110100100011101    1110100100011110    1110100100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59675 - 59679

  --1110100100100000    1110100100100001    1110100100100010    1110100100100011    1110100100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59680 - 59684

  --1110100100100101    1110100100100110    1110100100100111    1110100100101000    1110100100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59685 - 59689

  --1110100100101010    1110100100101011    1110100100101100    1110100100101101    1110100100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59690 - 59694

  --1110100100101111    1110100100110000    1110100100110001    1110100100110010    1110100100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59695 - 59699

  --1110100100110100    1110100100110101    1110100100110110    1110100100110111    1110100100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59700 - 59704

  --1110100100111001    1110100100111010    1110100100111011    1110100100111100    1110100100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59705 - 59709

  --1110100100111110    1110100100111111    1110100101000000    1110100101000001    1110100101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59710 - 59714

  --1110100101000011    1110100101000100    1110100101000101    1110100101000110    1110100101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59715 - 59719

  --1110100101001000    1110100101001001    1110100101001010    1110100101001011    1110100101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59720 - 59724

  --1110100101001101    1110100101001110    1110100101001111    1110100101010000    1110100101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59725 - 59729

  --1110100101010010    1110100101010011    1110100101010100    1110100101010101    1110100101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59730 - 59734

  --1110100101010111    1110100101011000    1110100101011001    1110100101011010    1110100101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59735 - 59739

  --1110100101011100    1110100101011101    1110100101011110    1110100101011111    1110100101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59740 - 59744

  --1110100101100001    1110100101100010    1110100101100011    1110100101100100    1110100101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59745 - 59749

  --1110100101100110    1110100101100111    1110100101101000    1110100101101001    1110100101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59750 - 59754

  --1110100101101011    1110100101101100    1110100101101101    1110100101101110    1110100101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59755 - 59759

  --1110100101110000    1110100101110001    1110100101110010    1110100101110011    1110100101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59760 - 59764

  --1110100101110101    1110100101110110    1110100101110111    1110100101111000    1110100101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59765 - 59769

  --1110100101111010    1110100101111011    1110100101111100    1110100101111101    1110100101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59770 - 59774

  --1110100101111111    1110100110000000    1110100110000001    1110100110000010    1110100110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59775 - 59779

  --1110100110000100    1110100110000101    1110100110000110    1110100110000111    1110100110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59780 - 59784

  --1110100110001001    1110100110001010    1110100110001011    1110100110001100    1110100110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59785 - 59789

  --1110100110001110    1110100110001111    1110100110010000    1110100110010001    1110100110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59790 - 59794

  --1110100110010011    1110100110010100    1110100110010101    1110100110010110    1110100110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59795 - 59799

  --1110100110011000    1110100110011001    1110100110011010    1110100110011011    1110100110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59800 - 59804

  --1110100110011101    1110100110011110    1110100110011111    1110100110100000    1110100110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59805 - 59809

  --1110100110100010    1110100110100011    1110100110100100    1110100110100101    1110100110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59810 - 59814

  --1110100110100111    1110100110101000    1110100110101001    1110100110101010    1110100110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59815 - 59819

  --1110100110101100    1110100110101101    1110100110101110    1110100110101111    1110100110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59820 - 59824

  --1110100110110001    1110100110110010    1110100110110011    1110100110110100    1110100110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59825 - 59829

  --1110100110110110    1110100110110111    1110100110111000    1110100110111001    1110100110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59830 - 59834

  --1110100110111011    1110100110111100    1110100110111101    1110100110111110    1110100110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59835 - 59839

  --1110100111000000    1110100111000001    1110100111000010    1110100111000011    1110100111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59840 - 59844

  --1110100111000101    1110100111000110    1110100111000111    1110100111001000    1110100111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59845 - 59849

  --1110100111001010    1110100111001011    1110100111001100    1110100111001101    1110100111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59850 - 59854

  --1110100111001111    1110100111010000    1110100111010001    1110100111010010    1110100111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59855 - 59859

  --1110100111010100    1110100111010101    1110100111010110    1110100111010111    1110100111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59860 - 59864

  --1110100111011001    1110100111011010    1110100111011011    1110100111011100    1110100111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59865 - 59869

  --1110100111011110    1110100111011111    1110100111100000    1110100111100001    1110100111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59870 - 59874

  --1110100111100011    1110100111100100    1110100111100101    1110100111100110    1110100111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59875 - 59879

  --1110100111101000    1110100111101001    1110100111101010    1110100111101011    1110100111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59880 - 59884

  --1110100111101101    1110100111101110    1110100111101111    1110100111110000    1110100111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59885 - 59889

  --1110100111110010    1110100111110011    1110100111110100    1110100111110101    1110100111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59890 - 59894

  --1110100111110111    1110100111111000    1110100111111001    1110100111111010    1110100111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59895 - 59899

  --1110100111111100    1110100111111101    1110100111111110    1110100111111111    1110101000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59900 - 59904

  --1110101000000001    1110101000000010    1110101000000011    1110101000000100    1110101000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59905 - 59909

  --1110101000000110    1110101000000111    1110101000001000    1110101000001001    1110101000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59910 - 59914

  --1110101000001011    1110101000001100    1110101000001101    1110101000001110    1110101000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59915 - 59919

  --1110101000010000    1110101000010001    1110101000010010    1110101000010011    1110101000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59920 - 59924

  --1110101000010101    1110101000010110    1110101000010111    1110101000011000    1110101000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59925 - 59929

  --1110101000011010    1110101000011011    1110101000011100    1110101000011101    1110101000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59930 - 59934

  --1110101000011111    1110101000100000    1110101000100001    1110101000100010    1110101000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59935 - 59939

  --1110101000100100    1110101000100101    1110101000100110    1110101000100111    1110101000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59940 - 59944

  --1110101000101001    1110101000101010    1110101000101011    1110101000101100    1110101000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59945 - 59949

  --1110101000101110    1110101000101111    1110101000110000    1110101000110001    1110101000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59950 - 59954

  --1110101000110011    1110101000110100    1110101000110101    1110101000110110    1110101000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59955 - 59959

  --1110101000111000    1110101000111001    1110101000111010    1110101000111011    1110101000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59960 - 59964

  --1110101000111101    1110101000111110    1110101000111111    1110101001000000    1110101001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59965 - 59969

  --1110101001000010    1110101001000011    1110101001000100    1110101001000101    1110101001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59970 - 59974

  --1110101001000111    1110101001001000    1110101001001001    1110101001001010    1110101001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59975 - 59979

  --1110101001001100    1110101001001101    1110101001001110    1110101001001111    1110101001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59980 - 59984

  --1110101001010001    1110101001010010    1110101001010011    1110101001010100    1110101001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59985 - 59989

  --1110101001010110    1110101001010111    1110101001011000    1110101001011001    1110101001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59990 - 59994

  --1110101001011011    1110101001011100    1110101001011101    1110101001011110    1110101001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 59995 - 59999

  --1110101001100000    1110101001100001    1110101001100010    1110101001100011    1110101001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60000 - 60004

  --1110101001100101    1110101001100110    1110101001100111    1110101001101000    1110101001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60005 - 60009

  --1110101001101010    1110101001101011    1110101001101100    1110101001101101    1110101001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60010 - 60014

  --1110101001101111    1110101001110000    1110101001110001    1110101001110010    1110101001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60015 - 60019

  --1110101001110100    1110101001110101    1110101001110110    1110101001110111    1110101001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60020 - 60024

  --1110101001111001    1110101001111010    1110101001111011    1110101001111100    1110101001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60025 - 60029

  --1110101001111110    1110101001111111    1110101010000000    1110101010000001    1110101010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60030 - 60034

  --1110101010000011    1110101010000100    1110101010000101    1110101010000110    1110101010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60035 - 60039

  --1110101010001000    1110101010001001    1110101010001010    1110101010001011    1110101010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60040 - 60044

  --1110101010001101    1110101010001110    1110101010001111    1110101010010000    1110101010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60045 - 60049

  --1110101010010010    1110101010010011    1110101010010100    1110101010010101    1110101010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60050 - 60054

  --1110101010010111    1110101010011000    1110101010011001    1110101010011010    1110101010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60055 - 60059

  --1110101010011100    1110101010011101    1110101010011110    1110101010011111    1110101010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60060 - 60064

  --1110101010100001    1110101010100010    1110101010100011    1110101010100100    1110101010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60065 - 60069

  --1110101010100110    1110101010100111    1110101010101000    1110101010101001    1110101010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60070 - 60074

  --1110101010101011    1110101010101100    1110101010101101    1110101010101110    1110101010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60075 - 60079

  --1110101010110000    1110101010110001    1110101010110010    1110101010110011    1110101010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60080 - 60084

  --1110101010110101    1110101010110110    1110101010110111    1110101010111000    1110101010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60085 - 60089

  --1110101010111010    1110101010111011    1110101010111100    1110101010111101    1110101010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60090 - 60094

  --1110101010111111    1110101011000000    1110101011000001    1110101011000010    1110101011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60095 - 60099

  --1110101011000100    1110101011000101    1110101011000110    1110101011000111    1110101011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60100 - 60104

  --1110101011001001    1110101011001010    1110101011001011    1110101011001100    1110101011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60105 - 60109

  --1110101011001110    1110101011001111    1110101011010000    1110101011010001    1110101011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60110 - 60114

  --1110101011010011    1110101011010100    1110101011010101    1110101011010110    1110101011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60115 - 60119

  --1110101011011000    1110101011011001    1110101011011010    1110101011011011    1110101011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60120 - 60124

  --1110101011011101    1110101011011110    1110101011011111    1110101011100000    1110101011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60125 - 60129

  --1110101011100010    1110101011100011    1110101011100100    1110101011100101    1110101011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60130 - 60134

  --1110101011100111    1110101011101000    1110101011101001    1110101011101010    1110101011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60135 - 60139

  --1110101011101100    1110101011101101    1110101011101110    1110101011101111    1110101011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60140 - 60144

  --1110101011110001    1110101011110010    1110101011110011    1110101011110100    1110101011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60145 - 60149

  --1110101011110110    1110101011110111    1110101011111000    1110101011111001    1110101011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60150 - 60154

  --1110101011111011    1110101011111100    1110101011111101    1110101011111110    1110101011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60155 - 60159

  --1110101100000000    1110101100000001    1110101100000010    1110101100000011    1110101100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60160 - 60164

  --1110101100000101    1110101100000110    1110101100000111    1110101100001000    1110101100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60165 - 60169

  --1110101100001010    1110101100001011    1110101100001100    1110101100001101    1110101100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60170 - 60174

  --1110101100001111    1110101100010000    1110101100010001    1110101100010010    1110101100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60175 - 60179

  --1110101100010100    1110101100010101    1110101100010110    1110101100010111    1110101100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60180 - 60184

  --1110101100011001    1110101100011010    1110101100011011    1110101100011100    1110101100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60185 - 60189

  --1110101100011110    1110101100011111    1110101100100000    1110101100100001    1110101100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60190 - 60194

  --1110101100100011    1110101100100100    1110101100100101    1110101100100110    1110101100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60195 - 60199

  --1110101100101000    1110101100101001    1110101100101010    1110101100101011    1110101100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60200 - 60204

  --1110101100101101    1110101100101110    1110101100101111    1110101100110000    1110101100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60205 - 60209

  --1110101100110010    1110101100110011    1110101100110100    1110101100110101    1110101100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60210 - 60214

  --1110101100110111    1110101100111000    1110101100111001    1110101100111010    1110101100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60215 - 60219

  --1110101100111100    1110101100111101    1110101100111110    1110101100111111    1110101101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60220 - 60224

  --1110101101000001    1110101101000010    1110101101000011    1110101101000100    1110101101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60225 - 60229

  --1110101101000110    1110101101000111    1110101101001000    1110101101001001    1110101101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60230 - 60234

  --1110101101001011    1110101101001100    1110101101001101    1110101101001110    1110101101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60235 - 60239

  --1110101101010000    1110101101010001    1110101101010010    1110101101010011    1110101101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60240 - 60244

  --1110101101010101    1110101101010110    1110101101010111    1110101101011000    1110101101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60245 - 60249

  --1110101101011010    1110101101011011    1110101101011100    1110101101011101    1110101101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60250 - 60254

  --1110101101011111    1110101101100000    1110101101100001    1110101101100010    1110101101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60255 - 60259

  --1110101101100100    1110101101100101    1110101101100110    1110101101100111    1110101101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60260 - 60264

  --1110101101101001    1110101101101010    1110101101101011    1110101101101100    1110101101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60265 - 60269

  --1110101101101110    1110101101101111    1110101101110000    1110101101110001    1110101101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60270 - 60274

  --1110101101110011    1110101101110100    1110101101110101    1110101101110110    1110101101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60275 - 60279

  --1110101101111000    1110101101111001    1110101101111010    1110101101111011    1110101101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60280 - 60284

  --1110101101111101    1110101101111110    1110101101111111    1110101110000000    1110101110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60285 - 60289

  --1110101110000010    1110101110000011    1110101110000100    1110101110000101    1110101110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60290 - 60294

  --1110101110000111    1110101110001000    1110101110001001    1110101110001010    1110101110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60295 - 60299

  --1110101110001100    1110101110001101    1110101110001110    1110101110001111    1110101110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60300 - 60304

  --1110101110010001    1110101110010010    1110101110010011    1110101110010100    1110101110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60305 - 60309

  --1110101110010110    1110101110010111    1110101110011000    1110101110011001    1110101110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60310 - 60314

  --1110101110011011    1110101110011100    1110101110011101    1110101110011110    1110101110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60315 - 60319

  --1110101110100000    1110101110100001    1110101110100010    1110101110100011    1110101110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60320 - 60324

  --1110101110100101    1110101110100110    1110101110100111    1110101110101000    1110101110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60325 - 60329

  --1110101110101010    1110101110101011    1110101110101100    1110101110101101    1110101110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60330 - 60334

  --1110101110101111    1110101110110000    1110101110110001    1110101110110010    1110101110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60335 - 60339

  --1110101110110100    1110101110110101    1110101110110110    1110101110110111    1110101110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60340 - 60344

  --1110101110111001    1110101110111010    1110101110111011    1110101110111100    1110101110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60345 - 60349

  --1110101110111110    1110101110111111    1110101111000000    1110101111000001    1110101111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60350 - 60354

  --1110101111000011    1110101111000100    1110101111000101    1110101111000110    1110101111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60355 - 60359

  --1110101111001000    1110101111001001    1110101111001010    1110101111001011    1110101111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60360 - 60364

  --1110101111001101    1110101111001110    1110101111001111    1110101111010000    1110101111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60365 - 60369

  --1110101111010010    1110101111010011    1110101111010100    1110101111010101    1110101111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60370 - 60374

  --1110101111010111    1110101111011000    1110101111011001    1110101111011010    1110101111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60375 - 60379

  --1110101111011100    1110101111011101    1110101111011110    1110101111011111    1110101111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60380 - 60384

  --1110101111100001    1110101111100010    1110101111100011    1110101111100100    1110101111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60385 - 60389

  --1110101111100110    1110101111100111    1110101111101000    1110101111101001    1110101111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60390 - 60394

  --1110101111101011    1110101111101100    1110101111101101    1110101111101110    1110101111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60395 - 60399

  --1110101111110000    1110101111110001    1110101111110010    1110101111110011    1110101111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60400 - 60404

  --1110101111110101    1110101111110110    1110101111110111    1110101111111000    1110101111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60405 - 60409

  --1110101111111010    1110101111111011    1110101111111100    1110101111111101    1110101111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60410 - 60414

  --1110101111111111    1110110000000000    1110110000000001    1110110000000010    1110110000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60415 - 60419

  --1110110000000100    1110110000000101    1110110000000110    1110110000000111    1110110000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60420 - 60424

  --1110110000001001    1110110000001010    1110110000001011    1110110000001100    1110110000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60425 - 60429

  --1110110000001110    1110110000001111    1110110000010000    1110110000010001    1110110000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60430 - 60434

  --1110110000010011    1110110000010100    1110110000010101    1110110000010110    1110110000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60435 - 60439

  --1110110000011000    1110110000011001    1110110000011010    1110110000011011    1110110000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60440 - 60444

  --1110110000011101    1110110000011110    1110110000011111    1110110000100000    1110110000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60445 - 60449

  --1110110000100010    1110110000100011    1110110000100100    1110110000100101    1110110000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60450 - 60454

  --1110110000100111    1110110000101000    1110110000101001    1110110000101010    1110110000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60455 - 60459

  --1110110000101100    1110110000101101    1110110000101110    1110110000101111    1110110000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60460 - 60464

  --1110110000110001    1110110000110010    1110110000110011    1110110000110100    1110110000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60465 - 60469

  --1110110000110110    1110110000110111    1110110000111000    1110110000111001    1110110000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60470 - 60474

  --1110110000111011    1110110000111100    1110110000111101    1110110000111110    1110110000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60475 - 60479

  --1110110001000000    1110110001000001    1110110001000010    1110110001000011    1110110001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60480 - 60484

  --1110110001000101    1110110001000110    1110110001000111    1110110001001000    1110110001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60485 - 60489

  --1110110001001010    1110110001001011    1110110001001100    1110110001001101    1110110001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60490 - 60494

  --1110110001001111    1110110001010000    1110110001010001    1110110001010010    1110110001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60495 - 60499

  --1110110001010100    1110110001010101    1110110001010110    1110110001010111    1110110001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60500 - 60504

  --1110110001011001    1110110001011010    1110110001011011    1110110001011100    1110110001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60505 - 60509

  --1110110001011110    1110110001011111    1110110001100000    1110110001100001    1110110001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60510 - 60514

  --1110110001100011    1110110001100100    1110110001100101    1110110001100110    1110110001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60515 - 60519

  --1110110001101000    1110110001101001    1110110001101010    1110110001101011    1110110001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60520 - 60524

  --1110110001101101    1110110001101110    1110110001101111    1110110001110000    1110110001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60525 - 60529

  --1110110001110010    1110110001110011    1110110001110100    1110110001110101    1110110001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60530 - 60534

  --1110110001110111    1110110001111000    1110110001111001    1110110001111010    1110110001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60535 - 60539

  --1110110001111100    1110110001111101    1110110001111110    1110110001111111    1110110010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60540 - 60544

  --1110110010000001    1110110010000010    1110110010000011    1110110010000100    1110110010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60545 - 60549

  --1110110010000110    1110110010000111    1110110010001000    1110110010001001    1110110010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60550 - 60554

  --1110110010001011    1110110010001100    1110110010001101    1110110010001110    1110110010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60555 - 60559

  --1110110010010000    1110110010010001    1110110010010010    1110110010010011    1110110010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60560 - 60564

  --1110110010010101    1110110010010110    1110110010010111    1110110010011000    1110110010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60565 - 60569

  --1110110010011010    1110110010011011    1110110010011100    1110110010011101    1110110010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60570 - 60574

  --1110110010011111    1110110010100000    1110110010100001    1110110010100010    1110110010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60575 - 60579

  --1110110010100100    1110110010100101    1110110010100110    1110110010100111    1110110010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60580 - 60584

  --1110110010101001    1110110010101010    1110110010101011    1110110010101100    1110110010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60585 - 60589

  --1110110010101110    1110110010101111    1110110010110000    1110110010110001    1110110010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60590 - 60594

  --1110110010110011    1110110010110100    1110110010110101    1110110010110110    1110110010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60595 - 60599

  --1110110010111000    1110110010111001    1110110010111010    1110110010111011    1110110010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60600 - 60604

  --1110110010111101    1110110010111110    1110110010111111    1110110011000000    1110110011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60605 - 60609

  --1110110011000010    1110110011000011    1110110011000100    1110110011000101    1110110011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60610 - 60614

  --1110110011000111    1110110011001000    1110110011001001    1110110011001010    1110110011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60615 - 60619

  --1110110011001100    1110110011001101    1110110011001110    1110110011001111    1110110011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60620 - 60624

  --1110110011010001    1110110011010010    1110110011010011    1110110011010100    1110110011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60625 - 60629

  --1110110011010110    1110110011010111    1110110011011000    1110110011011001    1110110011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60630 - 60634

  --1110110011011011    1110110011011100    1110110011011101    1110110011011110    1110110011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60635 - 60639

  --1110110011100000    1110110011100001    1110110011100010    1110110011100011    1110110011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60640 - 60644

  --1110110011100101    1110110011100110    1110110011100111    1110110011101000    1110110011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60645 - 60649

  --1110110011101010    1110110011101011    1110110011101100    1110110011101101    1110110011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60650 - 60654

  --1110110011101111    1110110011110000    1110110011110001    1110110011110010    1110110011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60655 - 60659

  --1110110011110100    1110110011110101    1110110011110110    1110110011110111    1110110011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60660 - 60664

  --1110110011111001    1110110011111010    1110110011111011    1110110011111100    1110110011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60665 - 60669

  --1110110011111110    1110110011111111    1110110100000000    1110110100000001    1110110100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60670 - 60674

  --1110110100000011    1110110100000100    1110110100000101    1110110100000110    1110110100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60675 - 60679

  --1110110100001000    1110110100001001    1110110100001010    1110110100001011    1110110100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60680 - 60684

  --1110110100001101    1110110100001110    1110110100001111    1110110100010000    1110110100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60685 - 60689

  --1110110100010010    1110110100010011    1110110100010100    1110110100010101    1110110100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60690 - 60694

  --1110110100010111    1110110100011000    1110110100011001    1110110100011010    1110110100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60695 - 60699

  --1110110100011100    1110110100011101    1110110100011110    1110110100011111    1110110100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60700 - 60704

  --1110110100100001    1110110100100010    1110110100100011    1110110100100100    1110110100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60705 - 60709

  --1110110100100110    1110110100100111    1110110100101000    1110110100101001    1110110100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60710 - 60714

  --1110110100101011    1110110100101100    1110110100101101    1110110100101110    1110110100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60715 - 60719

  --1110110100110000    1110110100110001    1110110100110010    1110110100110011    1110110100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60720 - 60724

  --1110110100110101    1110110100110110    1110110100110111    1110110100111000    1110110100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60725 - 60729

  --1110110100111010    1110110100111011    1110110100111100    1110110100111101    1110110100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60730 - 60734

  --1110110100111111    1110110101000000    1110110101000001    1110110101000010    1110110101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60735 - 60739

  --1110110101000100    1110110101000101    1110110101000110    1110110101000111    1110110101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60740 - 60744

  --1110110101001001    1110110101001010    1110110101001011    1110110101001100    1110110101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60745 - 60749

  --1110110101001110    1110110101001111    1110110101010000    1110110101010001    1110110101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60750 - 60754

  --1110110101010011    1110110101010100    1110110101010101    1110110101010110    1110110101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60755 - 60759

  --1110110101011000    1110110101011001    1110110101011010    1110110101011011    1110110101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60760 - 60764

  --1110110101011101    1110110101011110    1110110101011111    1110110101100000    1110110101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60765 - 60769

  --1110110101100010    1110110101100011    1110110101100100    1110110101100101    1110110101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60770 - 60774

  --1110110101100111    1110110101101000    1110110101101001    1110110101101010    1110110101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60775 - 60779

  --1110110101101100    1110110101101101    1110110101101110    1110110101101111    1110110101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60780 - 60784

  --1110110101110001    1110110101110010    1110110101110011    1110110101110100    1110110101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60785 - 60789

  --1110110101110110    1110110101110111    1110110101111000    1110110101111001    1110110101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60790 - 60794

  --1110110101111011    1110110101111100    1110110101111101    1110110101111110    1110110101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60795 - 60799

  --1110110110000000    1110110110000001    1110110110000010    1110110110000011    1110110110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60800 - 60804

  --1110110110000101    1110110110000110    1110110110000111    1110110110001000    1110110110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60805 - 60809

  --1110110110001010    1110110110001011    1110110110001100    1110110110001101    1110110110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60810 - 60814

  --1110110110001111    1110110110010000    1110110110010001    1110110110010010    1110110110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60815 - 60819

  --1110110110010100    1110110110010101    1110110110010110    1110110110010111    1110110110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60820 - 60824

  --1110110110011001    1110110110011010    1110110110011011    1110110110011100    1110110110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60825 - 60829

  --1110110110011110    1110110110011111    1110110110100000    1110110110100001    1110110110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60830 - 60834

  --1110110110100011    1110110110100100    1110110110100101    1110110110100110    1110110110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60835 - 60839

  --1110110110101000    1110110110101001    1110110110101010    1110110110101011    1110110110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60840 - 60844

  --1110110110101101    1110110110101110    1110110110101111    1110110110110000    1110110110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60845 - 60849

  --1110110110110010    1110110110110011    1110110110110100    1110110110110101    1110110110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60850 - 60854

  --1110110110110111    1110110110111000    1110110110111001    1110110110111010    1110110110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60855 - 60859

  --1110110110111100    1110110110111101    1110110110111110    1110110110111111    1110110111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60860 - 60864

  --1110110111000001    1110110111000010    1110110111000011    1110110111000100    1110110111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60865 - 60869

  --1110110111000110    1110110111000111    1110110111001000    1110110111001001    1110110111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60870 - 60874

  --1110110111001011    1110110111001100    1110110111001101    1110110111001110    1110110111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60875 - 60879

  --1110110111010000    1110110111010001    1110110111010010    1110110111010011    1110110111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60880 - 60884

  --1110110111010101    1110110111010110    1110110111010111    1110110111011000    1110110111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60885 - 60889

  --1110110111011010    1110110111011011    1110110111011100    1110110111011101    1110110111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60890 - 60894

  --1110110111011111    1110110111100000    1110110111100001    1110110111100010    1110110111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60895 - 60899

  --1110110111100100    1110110111100101    1110110111100110    1110110111100111    1110110111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60900 - 60904

  --1110110111101001    1110110111101010    1110110111101011    1110110111101100    1110110111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60905 - 60909

  --1110110111101110    1110110111101111    1110110111110000    1110110111110001    1110110111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60910 - 60914

  --1110110111110011    1110110111110100    1110110111110101    1110110111110110    1110110111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60915 - 60919

  --1110110111111000    1110110111111001    1110110111111010    1110110111111011    1110110111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60920 - 60924

  --1110110111111101    1110110111111110    1110110111111111    1110111000000000    1110111000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60925 - 60929

  --1110111000000010    1110111000000011    1110111000000100    1110111000000101    1110111000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60930 - 60934

  --1110111000000111    1110111000001000    1110111000001001    1110111000001010    1110111000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60935 - 60939

  --1110111000001100    1110111000001101    1110111000001110    1110111000001111    1110111000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60940 - 60944

  --1110111000010001    1110111000010010    1110111000010011    1110111000010100    1110111000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60945 - 60949

  --1110111000010110    1110111000010111    1110111000011000    1110111000011001    1110111000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60950 - 60954

  --1110111000011011    1110111000011100    1110111000011101    1110111000011110    1110111000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60955 - 60959

  --1110111000100000    1110111000100001    1110111000100010    1110111000100011    1110111000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60960 - 60964

  --1110111000100101    1110111000100110    1110111000100111    1110111000101000    1110111000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60965 - 60969

  --1110111000101010    1110111000101011    1110111000101100    1110111000101101    1110111000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60970 - 60974

  --1110111000101111    1110111000110000    1110111000110001    1110111000110010    1110111000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60975 - 60979

  --1110111000110100    1110111000110101    1110111000110110    1110111000110111    1110111000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60980 - 60984

  --1110111000111001    1110111000111010    1110111000111011    1110111000111100    1110111000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60985 - 60989

  --1110111000111110    1110111000111111    1110111001000000    1110111001000001    1110111001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60990 - 60994

  --1110111001000011    1110111001000100    1110111001000101    1110111001000110    1110111001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 60995 - 60999

  --1110111001001000    1110111001001001    1110111001001010    1110111001001011    1110111001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61000 - 61004

  --1110111001001101    1110111001001110    1110111001001111    1110111001010000    1110111001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61005 - 61009

  --1110111001010010    1110111001010011    1110111001010100    1110111001010101    1110111001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61010 - 61014

  --1110111001010111    1110111001011000    1110111001011001    1110111001011010    1110111001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61015 - 61019

  --1110111001011100    1110111001011101    1110111001011110    1110111001011111    1110111001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61020 - 61024

  --1110111001100001    1110111001100010    1110111001100011    1110111001100100    1110111001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61025 - 61029

  --1110111001100110    1110111001100111    1110111001101000    1110111001101001    1110111001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61030 - 61034

  --1110111001101011    1110111001101100    1110111001101101    1110111001101110    1110111001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61035 - 61039

  --1110111001110000    1110111001110001    1110111001110010    1110111001110011    1110111001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61040 - 61044

  --1110111001110101    1110111001110110    1110111001110111    1110111001111000    1110111001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61045 - 61049

  --1110111001111010    1110111001111011    1110111001111100    1110111001111101    1110111001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61050 - 61054

  --1110111001111111    1110111010000000    1110111010000001    1110111010000010    1110111010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61055 - 61059

  --1110111010000100    1110111010000101    1110111010000110    1110111010000111    1110111010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61060 - 61064

  --1110111010001001    1110111010001010    1110111010001011    1110111010001100    1110111010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61065 - 61069

  --1110111010001110    1110111010001111    1110111010010000    1110111010010001    1110111010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61070 - 61074

  --1110111010010011    1110111010010100    1110111010010101    1110111010010110    1110111010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61075 - 61079

  --1110111010011000    1110111010011001    1110111010011010    1110111010011011    1110111010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61080 - 61084

  --1110111010011101    1110111010011110    1110111010011111    1110111010100000    1110111010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61085 - 61089

  --1110111010100010    1110111010100011    1110111010100100    1110111010100101    1110111010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61090 - 61094

  --1110111010100111    1110111010101000    1110111010101001    1110111010101010    1110111010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61095 - 61099

  --1110111010101100    1110111010101101    1110111010101110    1110111010101111    1110111010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61100 - 61104

  --1110111010110001    1110111010110010    1110111010110011    1110111010110100    1110111010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61105 - 61109

  --1110111010110110    1110111010110111    1110111010111000    1110111010111001    1110111010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61110 - 61114

  --1110111010111011    1110111010111100    1110111010111101    1110111010111110    1110111010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61115 - 61119

  --1110111011000000    1110111011000001    1110111011000010    1110111011000011    1110111011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61120 - 61124

  --1110111011000101    1110111011000110    1110111011000111    1110111011001000    1110111011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61125 - 61129

  --1110111011001010    1110111011001011    1110111011001100    1110111011001101    1110111011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61130 - 61134

  --1110111011001111    1110111011010000    1110111011010001    1110111011010010    1110111011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61135 - 61139

  --1110111011010100    1110111011010101    1110111011010110    1110111011010111    1110111011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61140 - 61144

  --1110111011011001    1110111011011010    1110111011011011    1110111011011100    1110111011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61145 - 61149

  --1110111011011110    1110111011011111    1110111011100000    1110111011100001    1110111011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61150 - 61154

  --1110111011100011    1110111011100100    1110111011100101    1110111011100110    1110111011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61155 - 61159

  --1110111011101000    1110111011101001    1110111011101010    1110111011101011    1110111011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61160 - 61164

  --1110111011101101    1110111011101110    1110111011101111    1110111011110000    1110111011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61165 - 61169

  --1110111011110010    1110111011110011    1110111011110100    1110111011110101    1110111011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61170 - 61174

  --1110111011110111    1110111011111000    1110111011111001    1110111011111010    1110111011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61175 - 61179

  --1110111011111100    1110111011111101    1110111011111110    1110111011111111    1110111100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61180 - 61184

  --1110111100000001    1110111100000010    1110111100000011    1110111100000100    1110111100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61185 - 61189

  --1110111100000110    1110111100000111    1110111100001000    1110111100001001    1110111100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61190 - 61194

  --1110111100001011    1110111100001100    1110111100001101    1110111100001110    1110111100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61195 - 61199

  --1110111100010000    1110111100010001    1110111100010010    1110111100010011    1110111100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61200 - 61204

  --1110111100010101    1110111100010110    1110111100010111    1110111100011000    1110111100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61205 - 61209

  --1110111100011010    1110111100011011    1110111100011100    1110111100011101    1110111100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61210 - 61214

  --1110111100011111    1110111100100000    1110111100100001    1110111100100010    1110111100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61215 - 61219

  --1110111100100100    1110111100100101    1110111100100110    1110111100100111    1110111100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61220 - 61224

  --1110111100101001    1110111100101010    1110111100101011    1110111100101100    1110111100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61225 - 61229

  --1110111100101110    1110111100101111    1110111100110000    1110111100110001    1110111100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61230 - 61234

  --1110111100110011    1110111100110100    1110111100110101    1110111100110110    1110111100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61235 - 61239

  --1110111100111000    1110111100111001    1110111100111010    1110111100111011    1110111100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61240 - 61244

  --1110111100111101    1110111100111110    1110111100111111    1110111101000000    1110111101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61245 - 61249

  --1110111101000010    1110111101000011    1110111101000100    1110111101000101    1110111101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61250 - 61254

  --1110111101000111    1110111101001000    1110111101001001    1110111101001010    1110111101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61255 - 61259

  --1110111101001100    1110111101001101    1110111101001110    1110111101001111    1110111101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61260 - 61264

  --1110111101010001    1110111101010010    1110111101010011    1110111101010100    1110111101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61265 - 61269

  --1110111101010110    1110111101010111    1110111101011000    1110111101011001    1110111101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61270 - 61274

  --1110111101011011    1110111101011100    1110111101011101    1110111101011110    1110111101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61275 - 61279

  --1110111101100000    1110111101100001    1110111101100010    1110111101100011    1110111101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61280 - 61284

  --1110111101100101    1110111101100110    1110111101100111    1110111101101000    1110111101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61285 - 61289

  --1110111101101010    1110111101101011    1110111101101100    1110111101101101    1110111101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61290 - 61294

  --1110111101101111    1110111101110000    1110111101110001    1110111101110010    1110111101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61295 - 61299

  --1110111101110100    1110111101110101    1110111101110110    1110111101110111    1110111101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61300 - 61304

  --1110111101111001    1110111101111010    1110111101111011    1110111101111100    1110111101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61305 - 61309

  --1110111101111110    1110111101111111    1110111110000000    1110111110000001    1110111110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61310 - 61314

  --1110111110000011    1110111110000100    1110111110000101    1110111110000110    1110111110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61315 - 61319

  --1110111110001000    1110111110001001    1110111110001010    1110111110001011    1110111110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61320 - 61324

  --1110111110001101    1110111110001110    1110111110001111    1110111110010000    1110111110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61325 - 61329

  --1110111110010010    1110111110010011    1110111110010100    1110111110010101    1110111110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61330 - 61334

  --1110111110010111    1110111110011000    1110111110011001    1110111110011010    1110111110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61335 - 61339

  --1110111110011100    1110111110011101    1110111110011110    1110111110011111    1110111110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61340 - 61344

  --1110111110100001    1110111110100010    1110111110100011    1110111110100100    1110111110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61345 - 61349

  --1110111110100110    1110111110100111    1110111110101000    1110111110101001    1110111110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61350 - 61354

  --1110111110101011    1110111110101100    1110111110101101    1110111110101110    1110111110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61355 - 61359

  --1110111110110000    1110111110110001    1110111110110010    1110111110110011    1110111110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61360 - 61364

  --1110111110110101    1110111110110110    1110111110110111    1110111110111000    1110111110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61365 - 61369

  --1110111110111010    1110111110111011    1110111110111100    1110111110111101    1110111110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61370 - 61374

  --1110111110111111    1110111111000000    1110111111000001    1110111111000010    1110111111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61375 - 61379

  --1110111111000100    1110111111000101    1110111111000110    1110111111000111    1110111111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61380 - 61384

  --1110111111001001    1110111111001010    1110111111001011    1110111111001100    1110111111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61385 - 61389

  --1110111111001110    1110111111001111    1110111111010000    1110111111010001    1110111111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61390 - 61394

  --1110111111010011    1110111111010100    1110111111010101    1110111111010110    1110111111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61395 - 61399

  --1110111111011000    1110111111011001    1110111111011010    1110111111011011    1110111111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61400 - 61404

  --1110111111011101    1110111111011110    1110111111011111    1110111111100000    1110111111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61405 - 61409

  --1110111111100010    1110111111100011    1110111111100100    1110111111100101    1110111111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61410 - 61414

  --1110111111100111    1110111111101000    1110111111101001    1110111111101010    1110111111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61415 - 61419

  --1110111111101100    1110111111101101    1110111111101110    1110111111101111    1110111111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61420 - 61424

  --1110111111110001    1110111111110010    1110111111110011    1110111111110100    1110111111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61425 - 61429

  --1110111111110110    1110111111110111    1110111111111000    1110111111111001    1110111111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61430 - 61434

  --1110111111111011    1110111111111100    1110111111111101    1110111111111110    1110111111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61435 - 61439

  --1111000000000000    1111000000000001    1111000000000010    1111000000000011    1111000000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61440 - 61444

  --1111000000000101    1111000000000110    1111000000000111    1111000000001000    1111000000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61445 - 61449

  --1111000000001010    1111000000001011    1111000000001100    1111000000001101    1111000000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61450 - 61454

  --1111000000001111    1111000000010000    1111000000010001    1111000000010010    1111000000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61455 - 61459

  --1111000000010100    1111000000010101    1111000000010110    1111000000010111    1111000000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61460 - 61464

  --1111000000011001    1111000000011010    1111000000011011    1111000000011100    1111000000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61465 - 61469

  --1111000000011110    1111000000011111    1111000000100000    1111000000100001    1111000000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61470 - 61474

  --1111000000100011    1111000000100100    1111000000100101    1111000000100110    1111000000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61475 - 61479

  --1111000000101000    1111000000101001    1111000000101010    1111000000101011    1111000000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61480 - 61484

  --1111000000101101    1111000000101110    1111000000101111    1111000000110000    1111000000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61485 - 61489

  --1111000000110010    1111000000110011    1111000000110100    1111000000110101    1111000000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61490 - 61494

  --1111000000110111    1111000000111000    1111000000111001    1111000000111010    1111000000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61495 - 61499

  --1111000000111100    1111000000111101    1111000000111110    1111000000111111    1111000001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61500 - 61504

  --1111000001000001    1111000001000010    1111000001000011    1111000001000100    1111000001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61505 - 61509

  --1111000001000110    1111000001000111    1111000001001000    1111000001001001    1111000001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61510 - 61514

  --1111000001001011    1111000001001100    1111000001001101    1111000001001110    1111000001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61515 - 61519

  --1111000001010000    1111000001010001    1111000001010010    1111000001010011    1111000001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61520 - 61524

  --1111000001010101    1111000001010110    1111000001010111    1111000001011000    1111000001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61525 - 61529

  --1111000001011010    1111000001011011    1111000001011100    1111000001011101    1111000001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61530 - 61534

  --1111000001011111    1111000001100000    1111000001100001    1111000001100010    1111000001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61535 - 61539

  --1111000001100100    1111000001100101    1111000001100110    1111000001100111    1111000001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61540 - 61544

  --1111000001101001    1111000001101010    1111000001101011    1111000001101100    1111000001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61545 - 61549

  --1111000001101110    1111000001101111    1111000001110000    1111000001110001    1111000001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61550 - 61554

  --1111000001110011    1111000001110100    1111000001110101    1111000001110110    1111000001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61555 - 61559

  --1111000001111000    1111000001111001    1111000001111010    1111000001111011    1111000001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61560 - 61564

  --1111000001111101    1111000001111110    1111000001111111    1111000010000000    1111000010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61565 - 61569

  --1111000010000010    1111000010000011    1111000010000100    1111000010000101    1111000010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61570 - 61574

  --1111000010000111    1111000010001000    1111000010001001    1111000010001010    1111000010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61575 - 61579

  --1111000010001100    1111000010001101    1111000010001110    1111000010001111    1111000010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61580 - 61584

  --1111000010010001    1111000010010010    1111000010010011    1111000010010100    1111000010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61585 - 61589

  --1111000010010110    1111000010010111    1111000010011000    1111000010011001    1111000010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61590 - 61594

  --1111000010011011    1111000010011100    1111000010011101    1111000010011110    1111000010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61595 - 61599

  --1111000010100000    1111000010100001    1111000010100010    1111000010100011    1111000010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61600 - 61604

  --1111000010100101    1111000010100110    1111000010100111    1111000010101000    1111000010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61605 - 61609

  --1111000010101010    1111000010101011    1111000010101100    1111000010101101    1111000010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61610 - 61614

  --1111000010101111    1111000010110000    1111000010110001    1111000010110010    1111000010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61615 - 61619

  --1111000010110100    1111000010110101    1111000010110110    1111000010110111    1111000010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61620 - 61624

  --1111000010111001    1111000010111010    1111000010111011    1111000010111100    1111000010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61625 - 61629

  --1111000010111110    1111000010111111    1111000011000000    1111000011000001    1111000011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61630 - 61634

  --1111000011000011    1111000011000100    1111000011000101    1111000011000110    1111000011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61635 - 61639

  --1111000011001000    1111000011001001    1111000011001010    1111000011001011    1111000011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61640 - 61644

  --1111000011001101    1111000011001110    1111000011001111    1111000011010000    1111000011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61645 - 61649

  --1111000011010010    1111000011010011    1111000011010100    1111000011010101    1111000011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61650 - 61654

  --1111000011010111    1111000011011000    1111000011011001    1111000011011010    1111000011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61655 - 61659

  --1111000011011100    1111000011011101    1111000011011110    1111000011011111    1111000011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61660 - 61664

  --1111000011100001    1111000011100010    1111000011100011    1111000011100100    1111000011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61665 - 61669

  --1111000011100110    1111000011100111    1111000011101000    1111000011101001    1111000011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61670 - 61674

  --1111000011101011    1111000011101100    1111000011101101    1111000011101110    1111000011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61675 - 61679

  --1111000011110000    1111000011110001    1111000011110010    1111000011110011    1111000011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61680 - 61684

  --1111000011110101    1111000011110110    1111000011110111    1111000011111000    1111000011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61685 - 61689

  --1111000011111010    1111000011111011    1111000011111100    1111000011111101    1111000011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61690 - 61694

  --1111000011111111    1111000100000000    1111000100000001    1111000100000010    1111000100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61695 - 61699

  --1111000100000100    1111000100000101    1111000100000110    1111000100000111    1111000100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61700 - 61704

  --1111000100001001    1111000100001010    1111000100001011    1111000100001100    1111000100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61705 - 61709

  --1111000100001110    1111000100001111    1111000100010000    1111000100010001    1111000100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61710 - 61714

  --1111000100010011    1111000100010100    1111000100010101    1111000100010110    1111000100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61715 - 61719

  --1111000100011000    1111000100011001    1111000100011010    1111000100011011    1111000100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61720 - 61724

  --1111000100011101    1111000100011110    1111000100011111    1111000100100000    1111000100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61725 - 61729

  --1111000100100010    1111000100100011    1111000100100100    1111000100100101    1111000100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61730 - 61734

  --1111000100100111    1111000100101000    1111000100101001    1111000100101010    1111000100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61735 - 61739

  --1111000100101100    1111000100101101    1111000100101110    1111000100101111    1111000100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61740 - 61744

  --1111000100110001    1111000100110010    1111000100110011    1111000100110100    1111000100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61745 - 61749

  --1111000100110110    1111000100110111    1111000100111000    1111000100111001    1111000100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61750 - 61754

  --1111000100111011    1111000100111100    1111000100111101    1111000100111110    1111000100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61755 - 61759

  --1111000101000000    1111000101000001    1111000101000010    1111000101000011    1111000101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61760 - 61764

  --1111000101000101    1111000101000110    1111000101000111    1111000101001000    1111000101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61765 - 61769

  --1111000101001010    1111000101001011    1111000101001100    1111000101001101    1111000101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61770 - 61774

  --1111000101001111    1111000101010000    1111000101010001    1111000101010010    1111000101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61775 - 61779

  --1111000101010100    1111000101010101    1111000101010110    1111000101010111    1111000101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61780 - 61784

  --1111000101011001    1111000101011010    1111000101011011    1111000101011100    1111000101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61785 - 61789

  --1111000101011110    1111000101011111    1111000101100000    1111000101100001    1111000101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61790 - 61794

  --1111000101100011    1111000101100100    1111000101100101    1111000101100110    1111000101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61795 - 61799

  --1111000101101000    1111000101101001    1111000101101010    1111000101101011    1111000101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61800 - 61804

  --1111000101101101    1111000101101110    1111000101101111    1111000101110000    1111000101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61805 - 61809

  --1111000101110010    1111000101110011    1111000101110100    1111000101110101    1111000101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61810 - 61814

  --1111000101110111    1111000101111000    1111000101111001    1111000101111010    1111000101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61815 - 61819

  --1111000101111100    1111000101111101    1111000101111110    1111000101111111    1111000110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61820 - 61824

  --1111000110000001    1111000110000010    1111000110000011    1111000110000100    1111000110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61825 - 61829

  --1111000110000110    1111000110000111    1111000110001000    1111000110001001    1111000110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61830 - 61834

  --1111000110001011    1111000110001100    1111000110001101    1111000110001110    1111000110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61835 - 61839

  --1111000110010000    1111000110010001    1111000110010010    1111000110010011    1111000110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61840 - 61844

  --1111000110010101    1111000110010110    1111000110010111    1111000110011000    1111000110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61845 - 61849

  --1111000110011010    1111000110011011    1111000110011100    1111000110011101    1111000110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61850 - 61854

  --1111000110011111    1111000110100000    1111000110100001    1111000110100010    1111000110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61855 - 61859

  --1111000110100100    1111000110100101    1111000110100110    1111000110100111    1111000110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61860 - 61864

  --1111000110101001    1111000110101010    1111000110101011    1111000110101100    1111000110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61865 - 61869

  --1111000110101110    1111000110101111    1111000110110000    1111000110110001    1111000110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61870 - 61874

  --1111000110110011    1111000110110100    1111000110110101    1111000110110110    1111000110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61875 - 61879

  --1111000110111000    1111000110111001    1111000110111010    1111000110111011    1111000110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61880 - 61884

  --1111000110111101    1111000110111110    1111000110111111    1111000111000000    1111000111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61885 - 61889

  --1111000111000010    1111000111000011    1111000111000100    1111000111000101    1111000111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61890 - 61894

  --1111000111000111    1111000111001000    1111000111001001    1111000111001010    1111000111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61895 - 61899

  --1111000111001100    1111000111001101    1111000111001110    1111000111001111    1111000111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61900 - 61904

  --1111000111010001    1111000111010010    1111000111010011    1111000111010100    1111000111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61905 - 61909

  --1111000111010110    1111000111010111    1111000111011000    1111000111011001    1111000111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61910 - 61914

  --1111000111011011    1111000111011100    1111000111011101    1111000111011110    1111000111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61915 - 61919

  --1111000111100000    1111000111100001    1111000111100010    1111000111100011    1111000111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61920 - 61924

  --1111000111100101    1111000111100110    1111000111100111    1111000111101000    1111000111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61925 - 61929

  --1111000111101010    1111000111101011    1111000111101100    1111000111101101    1111000111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61930 - 61934

  --1111000111101111    1111000111110000    1111000111110001    1111000111110010    1111000111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61935 - 61939

  --1111000111110100    1111000111110101    1111000111110110    1111000111110111    1111000111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61940 - 61944

  --1111000111111001    1111000111111010    1111000111111011    1111000111111100    1111000111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61945 - 61949

  --1111000111111110    1111000111111111    1111001000000000    1111001000000001    1111001000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61950 - 61954

  --1111001000000011    1111001000000100    1111001000000101    1111001000000110    1111001000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61955 - 61959

  --1111001000001000    1111001000001001    1111001000001010    1111001000001011    1111001000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61960 - 61964

  --1111001000001101    1111001000001110    1111001000001111    1111001000010000    1111001000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61965 - 61969

  --1111001000010010    1111001000010011    1111001000010100    1111001000010101    1111001000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61970 - 61974

  --1111001000010111    1111001000011000    1111001000011001    1111001000011010    1111001000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61975 - 61979

  --1111001000011100    1111001000011101    1111001000011110    1111001000011111    1111001000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61980 - 61984

  --1111001000100001    1111001000100010    1111001000100011    1111001000100100    1111001000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61985 - 61989

  --1111001000100110    1111001000100111    1111001000101000    1111001000101001    1111001000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61990 - 61994

  --1111001000101011    1111001000101100    1111001000101101    1111001000101110    1111001000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 61995 - 61999

  --1111001000110000    1111001000110001    1111001000110010    1111001000110011    1111001000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62000 - 62004

  --1111001000110101    1111001000110110    1111001000110111    1111001000111000    1111001000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62005 - 62009

  --1111001000111010    1111001000111011    1111001000111100    1111001000111101    1111001000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62010 - 62014

  --1111001000111111    1111001001000000    1111001001000001    1111001001000010    1111001001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62015 - 62019

  --1111001001000100    1111001001000101    1111001001000110    1111001001000111    1111001001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62020 - 62024

  --1111001001001001    1111001001001010    1111001001001011    1111001001001100    1111001001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62025 - 62029

  --1111001001001110    1111001001001111    1111001001010000    1111001001010001    1111001001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62030 - 62034

  --1111001001010011    1111001001010100    1111001001010101    1111001001010110    1111001001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62035 - 62039

  --1111001001011000    1111001001011001    1111001001011010    1111001001011011    1111001001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62040 - 62044

  --1111001001011101    1111001001011110    1111001001011111    1111001001100000    1111001001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62045 - 62049

  --1111001001100010    1111001001100011    1111001001100100    1111001001100101    1111001001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62050 - 62054

  --1111001001100111    1111001001101000    1111001001101001    1111001001101010    1111001001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62055 - 62059

  --1111001001101100    1111001001101101    1111001001101110    1111001001101111    1111001001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62060 - 62064

  --1111001001110001    1111001001110010    1111001001110011    1111001001110100    1111001001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62065 - 62069

  --1111001001110110    1111001001110111    1111001001111000    1111001001111001    1111001001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62070 - 62074

  --1111001001111011    1111001001111100    1111001001111101    1111001001111110    1111001001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62075 - 62079

  --1111001010000000    1111001010000001    1111001010000010    1111001010000011    1111001010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62080 - 62084

  --1111001010000101    1111001010000110    1111001010000111    1111001010001000    1111001010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62085 - 62089

  --1111001010001010    1111001010001011    1111001010001100    1111001010001101    1111001010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62090 - 62094

  --1111001010001111    1111001010010000    1111001010010001    1111001010010010    1111001010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62095 - 62099

  --1111001010010100    1111001010010101    1111001010010110    1111001010010111    1111001010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62100 - 62104

  --1111001010011001    1111001010011010    1111001010011011    1111001010011100    1111001010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62105 - 62109

  --1111001010011110    1111001010011111    1111001010100000    1111001010100001    1111001010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62110 - 62114

  --1111001010100011    1111001010100100    1111001010100101    1111001010100110    1111001010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62115 - 62119

  --1111001010101000    1111001010101001    1111001010101010    1111001010101011    1111001010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62120 - 62124

  --1111001010101101    1111001010101110    1111001010101111    1111001010110000    1111001010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62125 - 62129

  --1111001010110010    1111001010110011    1111001010110100    1111001010110101    1111001010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62130 - 62134

  --1111001010110111    1111001010111000    1111001010111001    1111001010111010    1111001010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62135 - 62139

  --1111001010111100    1111001010111101    1111001010111110    1111001010111111    1111001011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62140 - 62144

  --1111001011000001    1111001011000010    1111001011000011    1111001011000100    1111001011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62145 - 62149

  --1111001011000110    1111001011000111    1111001011001000    1111001011001001    1111001011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62150 - 62154

  --1111001011001011    1111001011001100    1111001011001101    1111001011001110    1111001011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62155 - 62159

  --1111001011010000    1111001011010001    1111001011010010    1111001011010011    1111001011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62160 - 62164

  --1111001011010101    1111001011010110    1111001011010111    1111001011011000    1111001011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62165 - 62169

  --1111001011011010    1111001011011011    1111001011011100    1111001011011101    1111001011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62170 - 62174

  --1111001011011111    1111001011100000    1111001011100001    1111001011100010    1111001011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62175 - 62179

  --1111001011100100    1111001011100101    1111001011100110    1111001011100111    1111001011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62180 - 62184

  --1111001011101001    1111001011101010    1111001011101011    1111001011101100    1111001011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62185 - 62189

  --1111001011101110    1111001011101111    1111001011110000    1111001011110001    1111001011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62190 - 62194

  --1111001011110011    1111001011110100    1111001011110101    1111001011110110    1111001011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62195 - 62199

  --1111001011111000    1111001011111001    1111001011111010    1111001011111011    1111001011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62200 - 62204

  --1111001011111101    1111001011111110    1111001011111111    1111001100000000    1111001100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62205 - 62209

  --1111001100000010    1111001100000011    1111001100000100    1111001100000101    1111001100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62210 - 62214

  --1111001100000111    1111001100001000    1111001100001001    1111001100001010    1111001100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62215 - 62219

  --1111001100001100    1111001100001101    1111001100001110    1111001100001111    1111001100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62220 - 62224

  --1111001100010001    1111001100010010    1111001100010011    1111001100010100    1111001100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62225 - 62229

  --1111001100010110    1111001100010111    1111001100011000    1111001100011001    1111001100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62230 - 62234

  --1111001100011011    1111001100011100    1111001100011101    1111001100011110    1111001100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62235 - 62239

  --1111001100100000    1111001100100001    1111001100100010    1111001100100011    1111001100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62240 - 62244

  --1111001100100101    1111001100100110    1111001100100111    1111001100101000    1111001100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62245 - 62249

  --1111001100101010    1111001100101011    1111001100101100    1111001100101101    1111001100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62250 - 62254

  --1111001100101111    1111001100110000    1111001100110001    1111001100110010    1111001100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62255 - 62259

  --1111001100110100    1111001100110101    1111001100110110    1111001100110111    1111001100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62260 - 62264

  --1111001100111001    1111001100111010    1111001100111011    1111001100111100    1111001100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62265 - 62269

  --1111001100111110    1111001100111111    1111001101000000    1111001101000001    1111001101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62270 - 62274

  --1111001101000011    1111001101000100    1111001101000101    1111001101000110    1111001101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62275 - 62279

  --1111001101001000    1111001101001001    1111001101001010    1111001101001011    1111001101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62280 - 62284

  --1111001101001101    1111001101001110    1111001101001111    1111001101010000    1111001101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62285 - 62289

  --1111001101010010    1111001101010011    1111001101010100    1111001101010101    1111001101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62290 - 62294

  --1111001101010111    1111001101011000    1111001101011001    1111001101011010    1111001101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62295 - 62299

  --1111001101011100    1111001101011101    1111001101011110    1111001101011111    1111001101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62300 - 62304

  --1111001101100001    1111001101100010    1111001101100011    1111001101100100    1111001101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62305 - 62309

  --1111001101100110    1111001101100111    1111001101101000    1111001101101001    1111001101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62310 - 62314

  --1111001101101011    1111001101101100    1111001101101101    1111001101101110    1111001101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62315 - 62319

  --1111001101110000    1111001101110001    1111001101110010    1111001101110011    1111001101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62320 - 62324

  --1111001101110101    1111001101110110    1111001101110111    1111001101111000    1111001101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62325 - 62329

  --1111001101111010    1111001101111011    1111001101111100    1111001101111101    1111001101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62330 - 62334

  --1111001101111111    1111001110000000    1111001110000001    1111001110000010    1111001110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62335 - 62339

  --1111001110000100    1111001110000101    1111001110000110    1111001110000111    1111001110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62340 - 62344

  --1111001110001001    1111001110001010    1111001110001011    1111001110001100    1111001110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62345 - 62349

  --1111001110001110    1111001110001111    1111001110010000    1111001110010001    1111001110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62350 - 62354

  --1111001110010011    1111001110010100    1111001110010101    1111001110010110    1111001110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62355 - 62359

  --1111001110011000    1111001110011001    1111001110011010    1111001110011011    1111001110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62360 - 62364

  --1111001110011101    1111001110011110    1111001110011111    1111001110100000    1111001110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62365 - 62369

  --1111001110100010    1111001110100011    1111001110100100    1111001110100101    1111001110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62370 - 62374

  --1111001110100111    1111001110101000    1111001110101001    1111001110101010    1111001110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62375 - 62379

  --1111001110101100    1111001110101101    1111001110101110    1111001110101111    1111001110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62380 - 62384

  --1111001110110001    1111001110110010    1111001110110011    1111001110110100    1111001110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62385 - 62389

  --1111001110110110    1111001110110111    1111001110111000    1111001110111001    1111001110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62390 - 62394

  --1111001110111011    1111001110111100    1111001110111101    1111001110111110    1111001110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62395 - 62399

  --1111001111000000    1111001111000001    1111001111000010    1111001111000011    1111001111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62400 - 62404

  --1111001111000101    1111001111000110    1111001111000111    1111001111001000    1111001111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62405 - 62409

  --1111001111001010    1111001111001011    1111001111001100    1111001111001101    1111001111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62410 - 62414

  --1111001111001111    1111001111010000    1111001111010001    1111001111010010    1111001111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62415 - 62419

  --1111001111010100    1111001111010101    1111001111010110    1111001111010111    1111001111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62420 - 62424

  --1111001111011001    1111001111011010    1111001111011011    1111001111011100    1111001111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62425 - 62429

  --1111001111011110    1111001111011111    1111001111100000    1111001111100001    1111001111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62430 - 62434

  --1111001111100011    1111001111100100    1111001111100101    1111001111100110    1111001111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62435 - 62439

  --1111001111101000    1111001111101001    1111001111101010    1111001111101011    1111001111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62440 - 62444

  --1111001111101101    1111001111101110    1111001111101111    1111001111110000    1111001111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62445 - 62449

  --1111001111110010    1111001111110011    1111001111110100    1111001111110101    1111001111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62450 - 62454

  --1111001111110111    1111001111111000    1111001111111001    1111001111111010    1111001111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62455 - 62459

  --1111001111111100    1111001111111101    1111001111111110    1111001111111111    1111010000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62460 - 62464

  --1111010000000001    1111010000000010    1111010000000011    1111010000000100    1111010000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62465 - 62469

  --1111010000000110    1111010000000111    1111010000001000    1111010000001001    1111010000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62470 - 62474

  --1111010000001011    1111010000001100    1111010000001101    1111010000001110    1111010000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62475 - 62479

  --1111010000010000    1111010000010001    1111010000010010    1111010000010011    1111010000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62480 - 62484

  --1111010000010101    1111010000010110    1111010000010111    1111010000011000    1111010000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62485 - 62489

  --1111010000011010    1111010000011011    1111010000011100    1111010000011101    1111010000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62490 - 62494

  --1111010000011111    1111010000100000    1111010000100001    1111010000100010    1111010000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62495 - 62499

  --1111010000100100    1111010000100101    1111010000100110    1111010000100111    1111010000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62500 - 62504

  --1111010000101001    1111010000101010    1111010000101011    1111010000101100    1111010000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62505 - 62509

  --1111010000101110    1111010000101111    1111010000110000    1111010000110001    1111010000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62510 - 62514

  --1111010000110011    1111010000110100    1111010000110101    1111010000110110    1111010000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62515 - 62519

  --1111010000111000    1111010000111001    1111010000111010    1111010000111011    1111010000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62520 - 62524

  --1111010000111101    1111010000111110    1111010000111111    1111010001000000    1111010001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62525 - 62529

  --1111010001000010    1111010001000011    1111010001000100    1111010001000101    1111010001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62530 - 62534

  --1111010001000111    1111010001001000    1111010001001001    1111010001001010    1111010001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62535 - 62539

  --1111010001001100    1111010001001101    1111010001001110    1111010001001111    1111010001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62540 - 62544

  --1111010001010001    1111010001010010    1111010001010011    1111010001010100    1111010001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62545 - 62549

  --1111010001010110    1111010001010111    1111010001011000    1111010001011001    1111010001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62550 - 62554

  --1111010001011011    1111010001011100    1111010001011101    1111010001011110    1111010001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62555 - 62559

  --1111010001100000    1111010001100001    1111010001100010    1111010001100011    1111010001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62560 - 62564

  --1111010001100101    1111010001100110    1111010001100111    1111010001101000    1111010001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62565 - 62569

  --1111010001101010    1111010001101011    1111010001101100    1111010001101101    1111010001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62570 - 62574

  --1111010001101111    1111010001110000    1111010001110001    1111010001110010    1111010001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62575 - 62579

  --1111010001110100    1111010001110101    1111010001110110    1111010001110111    1111010001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62580 - 62584

  --1111010001111001    1111010001111010    1111010001111011    1111010001111100    1111010001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62585 - 62589

  --1111010001111110    1111010001111111    1111010010000000    1111010010000001    1111010010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62590 - 62594

  --1111010010000011    1111010010000100    1111010010000101    1111010010000110    1111010010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62595 - 62599

  --1111010010001000    1111010010001001    1111010010001010    1111010010001011    1111010010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62600 - 62604

  --1111010010001101    1111010010001110    1111010010001111    1111010010010000    1111010010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62605 - 62609

  --1111010010010010    1111010010010011    1111010010010100    1111010010010101    1111010010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62610 - 62614

  --1111010010010111    1111010010011000    1111010010011001    1111010010011010    1111010010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62615 - 62619

  --1111010010011100    1111010010011101    1111010010011110    1111010010011111    1111010010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62620 - 62624

  --1111010010100001    1111010010100010    1111010010100011    1111010010100100    1111010010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62625 - 62629

  --1111010010100110    1111010010100111    1111010010101000    1111010010101001    1111010010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62630 - 62634

  --1111010010101011    1111010010101100    1111010010101101    1111010010101110    1111010010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62635 - 62639

  --1111010010110000    1111010010110001    1111010010110010    1111010010110011    1111010010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62640 - 62644

  --1111010010110101    1111010010110110    1111010010110111    1111010010111000    1111010010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62645 - 62649

  --1111010010111010    1111010010111011    1111010010111100    1111010010111101    1111010010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62650 - 62654

  --1111010010111111    1111010011000000    1111010011000001    1111010011000010    1111010011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62655 - 62659

  --1111010011000100    1111010011000101    1111010011000110    1111010011000111    1111010011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62660 - 62664

  --1111010011001001    1111010011001010    1111010011001011    1111010011001100    1111010011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62665 - 62669

  --1111010011001110    1111010011001111    1111010011010000    1111010011010001    1111010011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62670 - 62674

  --1111010011010011    1111010011010100    1111010011010101    1111010011010110    1111010011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62675 - 62679

  --1111010011011000    1111010011011001    1111010011011010    1111010011011011    1111010011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62680 - 62684

  --1111010011011101    1111010011011110    1111010011011111    1111010011100000    1111010011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62685 - 62689

  --1111010011100010    1111010011100011    1111010011100100    1111010011100101    1111010011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62690 - 62694

  --1111010011100111    1111010011101000    1111010011101001    1111010011101010    1111010011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62695 - 62699

  --1111010011101100    1111010011101101    1111010011101110    1111010011101111    1111010011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62700 - 62704

  --1111010011110001    1111010011110010    1111010011110011    1111010011110100    1111010011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62705 - 62709

  --1111010011110110    1111010011110111    1111010011111000    1111010011111001    1111010011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62710 - 62714

  --1111010011111011    1111010011111100    1111010011111101    1111010011111110    1111010011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62715 - 62719

  --1111010100000000    1111010100000001    1111010100000010    1111010100000011    1111010100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62720 - 62724

  --1111010100000101    1111010100000110    1111010100000111    1111010100001000    1111010100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62725 - 62729

  --1111010100001010    1111010100001011    1111010100001100    1111010100001101    1111010100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62730 - 62734

  --1111010100001111    1111010100010000    1111010100010001    1111010100010010    1111010100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62735 - 62739

  --1111010100010100    1111010100010101    1111010100010110    1111010100010111    1111010100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62740 - 62744

  --1111010100011001    1111010100011010    1111010100011011    1111010100011100    1111010100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62745 - 62749

  --1111010100011110    1111010100011111    1111010100100000    1111010100100001    1111010100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62750 - 62754

  --1111010100100011    1111010100100100    1111010100100101    1111010100100110    1111010100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62755 - 62759

  --1111010100101000    1111010100101001    1111010100101010    1111010100101011    1111010100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62760 - 62764

  --1111010100101101    1111010100101110    1111010100101111    1111010100110000    1111010100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62765 - 62769

  --1111010100110010    1111010100110011    1111010100110100    1111010100110101    1111010100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62770 - 62774

  --1111010100110111    1111010100111000    1111010100111001    1111010100111010    1111010100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62775 - 62779

  --1111010100111100    1111010100111101    1111010100111110    1111010100111111    1111010101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62780 - 62784

  --1111010101000001    1111010101000010    1111010101000011    1111010101000100    1111010101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62785 - 62789

  --1111010101000110    1111010101000111    1111010101001000    1111010101001001    1111010101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62790 - 62794

  --1111010101001011    1111010101001100    1111010101001101    1111010101001110    1111010101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62795 - 62799

  --1111010101010000    1111010101010001    1111010101010010    1111010101010011    1111010101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62800 - 62804

  --1111010101010101    1111010101010110    1111010101010111    1111010101011000    1111010101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62805 - 62809

  --1111010101011010    1111010101011011    1111010101011100    1111010101011101    1111010101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62810 - 62814

  --1111010101011111    1111010101100000    1111010101100001    1111010101100010    1111010101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62815 - 62819

  --1111010101100100    1111010101100101    1111010101100110    1111010101100111    1111010101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62820 - 62824

  --1111010101101001    1111010101101010    1111010101101011    1111010101101100    1111010101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62825 - 62829

  --1111010101101110    1111010101101111    1111010101110000    1111010101110001    1111010101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62830 - 62834

  --1111010101110011    1111010101110100    1111010101110101    1111010101110110    1111010101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62835 - 62839

  --1111010101111000    1111010101111001    1111010101111010    1111010101111011    1111010101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62840 - 62844

  --1111010101111101    1111010101111110    1111010101111111    1111010110000000    1111010110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62845 - 62849

  --1111010110000010    1111010110000011    1111010110000100    1111010110000101    1111010110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62850 - 62854

  --1111010110000111    1111010110001000    1111010110001001    1111010110001010    1111010110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62855 - 62859

  --1111010110001100    1111010110001101    1111010110001110    1111010110001111    1111010110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62860 - 62864

  --1111010110010001    1111010110010010    1111010110010011    1111010110010100    1111010110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62865 - 62869

  --1111010110010110    1111010110010111    1111010110011000    1111010110011001    1111010110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62870 - 62874

  --1111010110011011    1111010110011100    1111010110011101    1111010110011110    1111010110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62875 - 62879

  --1111010110100000    1111010110100001    1111010110100010    1111010110100011    1111010110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62880 - 62884

  --1111010110100101    1111010110100110    1111010110100111    1111010110101000    1111010110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62885 - 62889

  --1111010110101010    1111010110101011    1111010110101100    1111010110101101    1111010110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62890 - 62894

  --1111010110101111    1111010110110000    1111010110110001    1111010110110010    1111010110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62895 - 62899

  --1111010110110100    1111010110110101    1111010110110110    1111010110110111    1111010110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62900 - 62904

  --1111010110111001    1111010110111010    1111010110111011    1111010110111100    1111010110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62905 - 62909

  --1111010110111110    1111010110111111    1111010111000000    1111010111000001    1111010111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62910 - 62914

  --1111010111000011    1111010111000100    1111010111000101    1111010111000110    1111010111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62915 - 62919

  --1111010111001000    1111010111001001    1111010111001010    1111010111001011    1111010111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62920 - 62924

  --1111010111001101    1111010111001110    1111010111001111    1111010111010000    1111010111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62925 - 62929

  --1111010111010010    1111010111010011    1111010111010100    1111010111010101    1111010111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62930 - 62934

  --1111010111010111    1111010111011000    1111010111011001    1111010111011010    1111010111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62935 - 62939

  --1111010111011100    1111010111011101    1111010111011110    1111010111011111    1111010111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62940 - 62944

  --1111010111100001    1111010111100010    1111010111100011    1111010111100100    1111010111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62945 - 62949

  --1111010111100110    1111010111100111    1111010111101000    1111010111101001    1111010111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62950 - 62954

  --1111010111101011    1111010111101100    1111010111101101    1111010111101110    1111010111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62955 - 62959

  --1111010111110000    1111010111110001    1111010111110010    1111010111110011    1111010111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62960 - 62964

  --1111010111110101    1111010111110110    1111010111110111    1111010111111000    1111010111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62965 - 62969

  --1111010111111010    1111010111111011    1111010111111100    1111010111111101    1111010111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62970 - 62974

  --1111010111111111    1111011000000000    1111011000000001    1111011000000010    1111011000000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62975 - 62979

  --1111011000000100    1111011000000101    1111011000000110    1111011000000111    1111011000001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62980 - 62984

  --1111011000001001    1111011000001010    1111011000001011    1111011000001100    1111011000001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62985 - 62989

  --1111011000001110    1111011000001111    1111011000010000    1111011000010001    1111011000010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62990 - 62994

  --1111011000010011    1111011000010100    1111011000010101    1111011000010110    1111011000010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 62995 - 62999

  --1111011000011000    1111011000011001    1111011000011010    1111011000011011    1111011000011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63000 - 63004

  --1111011000011101    1111011000011110    1111011000011111    1111011000100000    1111011000100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63005 - 63009

  --1111011000100010    1111011000100011    1111011000100100    1111011000100101    1111011000100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63010 - 63014

  --1111011000100111    1111011000101000    1111011000101001    1111011000101010    1111011000101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63015 - 63019

  --1111011000101100    1111011000101101    1111011000101110    1111011000101111    1111011000110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63020 - 63024

  --1111011000110001    1111011000110010    1111011000110011    1111011000110100    1111011000110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63025 - 63029

  --1111011000110110    1111011000110111    1111011000111000    1111011000111001    1111011000111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63030 - 63034

  --1111011000111011    1111011000111100    1111011000111101    1111011000111110    1111011000111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63035 - 63039

  --1111011001000000    1111011001000001    1111011001000010    1111011001000011    1111011001000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63040 - 63044

  --1111011001000101    1111011001000110    1111011001000111    1111011001001000    1111011001001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63045 - 63049

  --1111011001001010    1111011001001011    1111011001001100    1111011001001101    1111011001001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63050 - 63054

  --1111011001001111    1111011001010000    1111011001010001    1111011001010010    1111011001010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63055 - 63059

  --1111011001010100    1111011001010101    1111011001010110    1111011001010111    1111011001011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63060 - 63064

  --1111011001011001    1111011001011010    1111011001011011    1111011001011100    1111011001011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63065 - 63069

  --1111011001011110    1111011001011111    1111011001100000    1111011001100001    1111011001100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63070 - 63074

  --1111011001100011    1111011001100100    1111011001100101    1111011001100110    1111011001100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63075 - 63079

  --1111011001101000    1111011001101001    1111011001101010    1111011001101011    1111011001101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63080 - 63084

  --1111011001101101    1111011001101110    1111011001101111    1111011001110000    1111011001110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63085 - 63089

  --1111011001110010    1111011001110011    1111011001110100    1111011001110101    1111011001110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63090 - 63094

  --1111011001110111    1111011001111000    1111011001111001    1111011001111010    1111011001111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63095 - 63099

  --1111011001111100    1111011001111101    1111011001111110    1111011001111111    1111011010000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63100 - 63104

  --1111011010000001    1111011010000010    1111011010000011    1111011010000100    1111011010000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63105 - 63109

  --1111011010000110    1111011010000111    1111011010001000    1111011010001001    1111011010001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63110 - 63114

  --1111011010001011    1111011010001100    1111011010001101    1111011010001110    1111011010001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63115 - 63119

  --1111011010010000    1111011010010001    1111011010010010    1111011010010011    1111011010010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63120 - 63124

  --1111011010010101    1111011010010110    1111011010010111    1111011010011000    1111011010011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63125 - 63129

  --1111011010011010    1111011010011011    1111011010011100    1111011010011101    1111011010011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63130 - 63134

  --1111011010011111    1111011010100000    1111011010100001    1111011010100010    1111011010100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63135 - 63139

  --1111011010100100    1111011010100101    1111011010100110    1111011010100111    1111011010101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63140 - 63144

  --1111011010101001    1111011010101010    1111011010101011    1111011010101100    1111011010101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63145 - 63149

  --1111011010101110    1111011010101111    1111011010110000    1111011010110001    1111011010110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63150 - 63154

  --1111011010110011    1111011010110100    1111011010110101    1111011010110110    1111011010110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63155 - 63159

  --1111011010111000    1111011010111001    1111011010111010    1111011010111011    1111011010111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63160 - 63164

  --1111011010111101    1111011010111110    1111011010111111    1111011011000000    1111011011000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63165 - 63169

  --1111011011000010    1111011011000011    1111011011000100    1111011011000101    1111011011000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63170 - 63174

  --1111011011000111    1111011011001000    1111011011001001    1111011011001010    1111011011001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63175 - 63179

  --1111011011001100    1111011011001101    1111011011001110    1111011011001111    1111011011010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63180 - 63184

  --1111011011010001    1111011011010010    1111011011010011    1111011011010100    1111011011010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63185 - 63189

  --1111011011010110    1111011011010111    1111011011011000    1111011011011001    1111011011011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63190 - 63194

  --1111011011011011    1111011011011100    1111011011011101    1111011011011110    1111011011011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63195 - 63199

  --1111011011100000    1111011011100001    1111011011100010    1111011011100011    1111011011100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63200 - 63204

  --1111011011100101    1111011011100110    1111011011100111    1111011011101000    1111011011101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63205 - 63209

  --1111011011101010    1111011011101011    1111011011101100    1111011011101101    1111011011101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63210 - 63214

  --1111011011101111    1111011011110000    1111011011110001    1111011011110010    1111011011110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63215 - 63219

  --1111011011110100    1111011011110101    1111011011110110    1111011011110111    1111011011111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63220 - 63224

  --1111011011111001    1111011011111010    1111011011111011    1111011011111100    1111011011111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63225 - 63229

  --1111011011111110    1111011011111111    1111011100000000    1111011100000001    1111011100000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63230 - 63234

  --1111011100000011    1111011100000100    1111011100000101    1111011100000110    1111011100000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63235 - 63239

  --1111011100001000    1111011100001001    1111011100001010    1111011100001011    1111011100001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63240 - 63244

  --1111011100001101    1111011100001110    1111011100001111    1111011100010000    1111011100010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63245 - 63249

  --1111011100010010    1111011100010011    1111011100010100    1111011100010101    1111011100010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63250 - 63254

  --1111011100010111    1111011100011000    1111011100011001    1111011100011010    1111011100011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63255 - 63259

  --1111011100011100    1111011100011101    1111011100011110    1111011100011111    1111011100100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63260 - 63264

  --1111011100100001    1111011100100010    1111011100100011    1111011100100100    1111011100100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63265 - 63269

  --1111011100100110    1111011100100111    1111011100101000    1111011100101001    1111011100101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63270 - 63274

  --1111011100101011    1111011100101100    1111011100101101    1111011100101110    1111011100101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63275 - 63279

  --1111011100110000    1111011100110001    1111011100110010    1111011100110011    1111011100110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63280 - 63284

  --1111011100110101    1111011100110110    1111011100110111    1111011100111000    1111011100111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63285 - 63289

  --1111011100111010    1111011100111011    1111011100111100    1111011100111101    1111011100111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63290 - 63294

  --1111011100111111    1111011101000000    1111011101000001    1111011101000010    1111011101000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63295 - 63299

  --1111011101000100    1111011101000101    1111011101000110    1111011101000111    1111011101001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63300 - 63304

  --1111011101001001    1111011101001010    1111011101001011    1111011101001100    1111011101001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63305 - 63309

  --1111011101001110    1111011101001111    1111011101010000    1111011101010001    1111011101010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63310 - 63314

  --1111011101010011    1111011101010100    1111011101010101    1111011101010110    1111011101010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63315 - 63319

  --1111011101011000    1111011101011001    1111011101011010    1111011101011011    1111011101011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63320 - 63324

  --1111011101011101    1111011101011110    1111011101011111    1111011101100000    1111011101100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63325 - 63329

  --1111011101100010    1111011101100011    1111011101100100    1111011101100101    1111011101100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63330 - 63334

  --1111011101100111    1111011101101000    1111011101101001    1111011101101010    1111011101101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63335 - 63339

  --1111011101101100    1111011101101101    1111011101101110    1111011101101111    1111011101110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63340 - 63344

  --1111011101110001    1111011101110010    1111011101110011    1111011101110100    1111011101110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63345 - 63349

  --1111011101110110    1111011101110111    1111011101111000    1111011101111001    1111011101111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63350 - 63354

  --1111011101111011    1111011101111100    1111011101111101    1111011101111110    1111011101111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63355 - 63359

  --1111011110000000    1111011110000001    1111011110000010    1111011110000011    1111011110000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63360 - 63364

  --1111011110000101    1111011110000110    1111011110000111    1111011110001000    1111011110001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63365 - 63369

  --1111011110001010    1111011110001011    1111011110001100    1111011110001101    1111011110001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63370 - 63374

  --1111011110001111    1111011110010000    1111011110010001    1111011110010010    1111011110010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63375 - 63379

  --1111011110010100    1111011110010101    1111011110010110    1111011110010111    1111011110011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63380 - 63384

  --1111011110011001    1111011110011010    1111011110011011    1111011110011100    1111011110011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63385 - 63389

  --1111011110011110    1111011110011111    1111011110100000    1111011110100001    1111011110100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63390 - 63394

  --1111011110100011    1111011110100100    1111011110100101    1111011110100110    1111011110100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63395 - 63399

  --1111011110101000    1111011110101001    1111011110101010    1111011110101011    1111011110101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63400 - 63404

  --1111011110101101    1111011110101110    1111011110101111    1111011110110000    1111011110110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63405 - 63409

  --1111011110110010    1111011110110011    1111011110110100    1111011110110101    1111011110110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63410 - 63414

  --1111011110110111    1111011110111000    1111011110111001    1111011110111010    1111011110111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63415 - 63419

  --1111011110111100    1111011110111101    1111011110111110    1111011110111111    1111011111000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63420 - 63424

  --1111011111000001    1111011111000010    1111011111000011    1111011111000100    1111011111000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63425 - 63429

  --1111011111000110    1111011111000111    1111011111001000    1111011111001001    1111011111001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63430 - 63434

  --1111011111001011    1111011111001100    1111011111001101    1111011111001110    1111011111001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63435 - 63439

  --1111011111010000    1111011111010001    1111011111010010    1111011111010011    1111011111010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63440 - 63444

  --1111011111010101    1111011111010110    1111011111010111    1111011111011000    1111011111011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63445 - 63449

  --1111011111011010    1111011111011011    1111011111011100    1111011111011101    1111011111011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63450 - 63454

  --1111011111011111    1111011111100000    1111011111100001    1111011111100010    1111011111100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63455 - 63459

  --1111011111100100    1111011111100101    1111011111100110    1111011111100111    1111011111101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63460 - 63464

  --1111011111101001    1111011111101010    1111011111101011    1111011111101100    1111011111101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63465 - 63469

  --1111011111101110    1111011111101111    1111011111110000    1111011111110001    1111011111110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63470 - 63474

  --1111011111110011    1111011111110100    1111011111110101    1111011111110110    1111011111110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63475 - 63479

  --1111011111111000    1111011111111001    1111011111111010    1111011111111011    1111011111111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63480 - 63484

  --1111011111111101    1111011111111110    1111011111111111    1111100000000000    1111100000000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63485 - 63489

  --1111100000000010    1111100000000011    1111100000000100    1111100000000101    1111100000000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63490 - 63494

  --1111100000000111    1111100000001000    1111100000001001    1111100000001010    1111100000001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63495 - 63499

  --1111100000001100    1111100000001101    1111100000001110    1111100000001111    1111100000010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63500 - 63504

  --1111100000010001    1111100000010010    1111100000010011    1111100000010100    1111100000010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63505 - 63509

  --1111100000010110    1111100000010111    1111100000011000    1111100000011001    1111100000011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63510 - 63514

  --1111100000011011    1111100000011100    1111100000011101    1111100000011110    1111100000011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63515 - 63519

  --1111100000100000    1111100000100001    1111100000100010    1111100000100011    1111100000100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63520 - 63524

  --1111100000100101    1111100000100110    1111100000100111    1111100000101000    1111100000101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63525 - 63529

  --1111100000101010    1111100000101011    1111100000101100    1111100000101101    1111100000101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63530 - 63534

  --1111100000101111    1111100000110000    1111100000110001    1111100000110010    1111100000110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63535 - 63539

  --1111100000110100    1111100000110101    1111100000110110    1111100000110111    1111100000111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63540 - 63544

  --1111100000111001    1111100000111010    1111100000111011    1111100000111100    1111100000111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63545 - 63549

  --1111100000111110    1111100000111111    1111100001000000    1111100001000001    1111100001000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63550 - 63554

  --1111100001000011    1111100001000100    1111100001000101    1111100001000110    1111100001000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63555 - 63559

  --1111100001001000    1111100001001001    1111100001001010    1111100001001011    1111100001001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63560 - 63564

  --1111100001001101    1111100001001110    1111100001001111    1111100001010000    1111100001010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63565 - 63569

  --1111100001010010    1111100001010011    1111100001010100    1111100001010101    1111100001010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63570 - 63574

  --1111100001010111    1111100001011000    1111100001011001    1111100001011010    1111100001011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63575 - 63579

  --1111100001011100    1111100001011101    1111100001011110    1111100001011111    1111100001100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63580 - 63584

  --1111100001100001    1111100001100010    1111100001100011    1111100001100100    1111100001100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63585 - 63589

  --1111100001100110    1111100001100111    1111100001101000    1111100001101001    1111100001101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63590 - 63594

  --1111100001101011    1111100001101100    1111100001101101    1111100001101110    1111100001101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63595 - 63599

  --1111100001110000    1111100001110001    1111100001110010    1111100001110011    1111100001110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63600 - 63604

  --1111100001110101    1111100001110110    1111100001110111    1111100001111000    1111100001111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63605 - 63609

  --1111100001111010    1111100001111011    1111100001111100    1111100001111101    1111100001111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63610 - 63614

  --1111100001111111    1111100010000000    1111100010000001    1111100010000010    1111100010000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63615 - 63619

  --1111100010000100    1111100010000101    1111100010000110    1111100010000111    1111100010001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63620 - 63624

  --1111100010001001    1111100010001010    1111100010001011    1111100010001100    1111100010001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63625 - 63629

  --1111100010001110    1111100010001111    1111100010010000    1111100010010001    1111100010010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63630 - 63634

  --1111100010010011    1111100010010100    1111100010010101    1111100010010110    1111100010010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63635 - 63639

  --1111100010011000    1111100010011001    1111100010011010    1111100010011011    1111100010011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63640 - 63644

  --1111100010011101    1111100010011110    1111100010011111    1111100010100000    1111100010100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63645 - 63649

  --1111100010100010    1111100010100011    1111100010100100    1111100010100101    1111100010100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63650 - 63654

  --1111100010100111    1111100010101000    1111100010101001    1111100010101010    1111100010101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63655 - 63659

  --1111100010101100    1111100010101101    1111100010101110    1111100010101111    1111100010110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63660 - 63664

  --1111100010110001    1111100010110010    1111100010110011    1111100010110100    1111100010110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63665 - 63669

  --1111100010110110    1111100010110111    1111100010111000    1111100010111001    1111100010111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63670 - 63674

  --1111100010111011    1111100010111100    1111100010111101    1111100010111110    1111100010111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63675 - 63679

  --1111100011000000    1111100011000001    1111100011000010    1111100011000011    1111100011000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63680 - 63684

  --1111100011000101    1111100011000110    1111100011000111    1111100011001000    1111100011001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63685 - 63689

  --1111100011001010    1111100011001011    1111100011001100    1111100011001101    1111100011001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63690 - 63694

  --1111100011001111    1111100011010000    1111100011010001    1111100011010010    1111100011010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63695 - 63699

  --1111100011010100    1111100011010101    1111100011010110    1111100011010111    1111100011011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63700 - 63704

  --1111100011011001    1111100011011010    1111100011011011    1111100011011100    1111100011011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63705 - 63709

  --1111100011011110    1111100011011111    1111100011100000    1111100011100001    1111100011100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63710 - 63714

  --1111100011100011    1111100011100100    1111100011100101    1111100011100110    1111100011100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63715 - 63719

  --1111100011101000    1111100011101001    1111100011101010    1111100011101011    1111100011101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63720 - 63724

  --1111100011101101    1111100011101110    1111100011101111    1111100011110000    1111100011110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63725 - 63729

  --1111100011110010    1111100011110011    1111100011110100    1111100011110101    1111100011110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63730 - 63734

  --1111100011110111    1111100011111000    1111100011111001    1111100011111010    1111100011111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63735 - 63739

  --1111100011111100    1111100011111101    1111100011111110    1111100011111111    1111100100000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63740 - 63744

  --1111100100000001    1111100100000010    1111100100000011    1111100100000100    1111100100000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63745 - 63749

  --1111100100000110    1111100100000111    1111100100001000    1111100100001001    1111100100001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63750 - 63754

  --1111100100001011    1111100100001100    1111100100001101    1111100100001110    1111100100001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63755 - 63759

  --1111100100010000    1111100100010001    1111100100010010    1111100100010011    1111100100010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63760 - 63764

  --1111100100010101    1111100100010110    1111100100010111    1111100100011000    1111100100011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63765 - 63769

  --1111100100011010    1111100100011011    1111100100011100    1111100100011101    1111100100011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63770 - 63774

  --1111100100011111    1111100100100000    1111100100100001    1111100100100010    1111100100100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63775 - 63779

  --1111100100100100    1111100100100101    1111100100100110    1111100100100111    1111100100101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63780 - 63784

  --1111100100101001    1111100100101010    1111100100101011    1111100100101100    1111100100101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63785 - 63789

  --1111100100101110    1111100100101111    1111100100110000    1111100100110001    1111100100110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63790 - 63794

  --1111100100110011    1111100100110100    1111100100110101    1111100100110110    1111100100110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63795 - 63799

  --1111100100111000    1111100100111001    1111100100111010    1111100100111011    1111100100111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63800 - 63804

  --1111100100111101    1111100100111110    1111100100111111    1111100101000000    1111100101000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63805 - 63809

  --1111100101000010    1111100101000011    1111100101000100    1111100101000101    1111100101000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63810 - 63814

  --1111100101000111    1111100101001000    1111100101001001    1111100101001010    1111100101001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63815 - 63819

  --1111100101001100    1111100101001101    1111100101001110    1111100101001111    1111100101010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63820 - 63824

  --1111100101010001    1111100101010010    1111100101010011    1111100101010100    1111100101010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63825 - 63829

  --1111100101010110    1111100101010111    1111100101011000    1111100101011001    1111100101011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63830 - 63834

  --1111100101011011    1111100101011100    1111100101011101    1111100101011110    1111100101011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63835 - 63839

  --1111100101100000    1111100101100001    1111100101100010    1111100101100011    1111100101100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63840 - 63844

  --1111100101100101    1111100101100110    1111100101100111    1111100101101000    1111100101101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63845 - 63849

  --1111100101101010    1111100101101011    1111100101101100    1111100101101101    1111100101101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63850 - 63854

  --1111100101101111    1111100101110000    1111100101110001    1111100101110010    1111100101110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63855 - 63859

  --1111100101110100    1111100101110101    1111100101110110    1111100101110111    1111100101111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63860 - 63864

  --1111100101111001    1111100101111010    1111100101111011    1111100101111100    1111100101111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63865 - 63869

  --1111100101111110    1111100101111111    1111100110000000    1111100110000001    1111100110000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63870 - 63874

  --1111100110000011    1111100110000100    1111100110000101    1111100110000110    1111100110000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63875 - 63879

  --1111100110001000    1111100110001001    1111100110001010    1111100110001011    1111100110001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63880 - 63884

  --1111100110001101    1111100110001110    1111100110001111    1111100110010000    1111100110010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63885 - 63889

  --1111100110010010    1111100110010011    1111100110010100    1111100110010101    1111100110010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63890 - 63894

  --1111100110010111    1111100110011000    1111100110011001    1111100110011010    1111100110011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63895 - 63899

  --1111100110011100    1111100110011101    1111100110011110    1111100110011111    1111100110100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63900 - 63904

  --1111100110100001    1111100110100010    1111100110100011    1111100110100100    1111100110100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63905 - 63909

  --1111100110100110    1111100110100111    1111100110101000    1111100110101001    1111100110101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63910 - 63914

  --1111100110101011    1111100110101100    1111100110101101    1111100110101110    1111100110101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63915 - 63919

  --1111100110110000    1111100110110001    1111100110110010    1111100110110011    1111100110110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63920 - 63924

  --1111100110110101    1111100110110110    1111100110110111    1111100110111000    1111100110111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63925 - 63929

  --1111100110111010    1111100110111011    1111100110111100    1111100110111101    1111100110111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63930 - 63934

  --1111100110111111    1111100111000000    1111100111000001    1111100111000010    1111100111000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63935 - 63939

  --1111100111000100    1111100111000101    1111100111000110    1111100111000111    1111100111001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63940 - 63944

  --1111100111001001    1111100111001010    1111100111001011    1111100111001100    1111100111001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63945 - 63949

  --1111100111001110    1111100111001111    1111100111010000    1111100111010001    1111100111010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63950 - 63954

  --1111100111010011    1111100111010100    1111100111010101    1111100111010110    1111100111010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63955 - 63959

  --1111100111011000    1111100111011001    1111100111011010    1111100111011011    1111100111011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63960 - 63964

  --1111100111011101    1111100111011110    1111100111011111    1111100111100000    1111100111100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63965 - 63969

  --1111100111100010    1111100111100011    1111100111100100    1111100111100101    1111100111100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63970 - 63974

  --1111100111100111    1111100111101000    1111100111101001    1111100111101010    1111100111101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63975 - 63979

  --1111100111101100    1111100111101101    1111100111101110    1111100111101111    1111100111110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63980 - 63984

  --1111100111110001    1111100111110010    1111100111110011    1111100111110100    1111100111110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63985 - 63989

  --1111100111110110    1111100111110111    1111100111111000    1111100111111001    1111100111111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63990 - 63994

  --1111100111111011    1111100111111100    1111100111111101    1111100111111110    1111100111111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 63995 - 63999

  --1111101000000000    1111101000000001    1111101000000010    1111101000000011    1111101000000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64000 - 64004

  --1111101000000101    1111101000000110    1111101000000111    1111101000001000    1111101000001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64005 - 64009

  --1111101000001010    1111101000001011    1111101000001100    1111101000001101    1111101000001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64010 - 64014

  --1111101000001111    1111101000010000    1111101000010001    1111101000010010    1111101000010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64015 - 64019

  --1111101000010100    1111101000010101    1111101000010110    1111101000010111    1111101000011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64020 - 64024

  --1111101000011001    1111101000011010    1111101000011011    1111101000011100    1111101000011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64025 - 64029

  --1111101000011110    1111101000011111    1111101000100000    1111101000100001    1111101000100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64030 - 64034

  --1111101000100011    1111101000100100    1111101000100101    1111101000100110    1111101000100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64035 - 64039

  --1111101000101000    1111101000101001    1111101000101010    1111101000101011    1111101000101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64040 - 64044

  --1111101000101101    1111101000101110    1111101000101111    1111101000110000    1111101000110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64045 - 64049

  --1111101000110010    1111101000110011    1111101000110100    1111101000110101    1111101000110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64050 - 64054

  --1111101000110111    1111101000111000    1111101000111001    1111101000111010    1111101000111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64055 - 64059

  --1111101000111100    1111101000111101    1111101000111110    1111101000111111    1111101001000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64060 - 64064

  --1111101001000001    1111101001000010    1111101001000011    1111101001000100    1111101001000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64065 - 64069

  --1111101001000110    1111101001000111    1111101001001000    1111101001001001    1111101001001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64070 - 64074

  --1111101001001011    1111101001001100    1111101001001101    1111101001001110    1111101001001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64075 - 64079

  --1111101001010000    1111101001010001    1111101001010010    1111101001010011    1111101001010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64080 - 64084

  --1111101001010101    1111101001010110    1111101001010111    1111101001011000    1111101001011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64085 - 64089

  --1111101001011010    1111101001011011    1111101001011100    1111101001011101    1111101001011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64090 - 64094

  --1111101001011111    1111101001100000    1111101001100001    1111101001100010    1111101001100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64095 - 64099

  --1111101001100100    1111101001100101    1111101001100110    1111101001100111    1111101001101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64100 - 64104

  --1111101001101001    1111101001101010    1111101001101011    1111101001101100    1111101001101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64105 - 64109

  --1111101001101110    1111101001101111    1111101001110000    1111101001110001    1111101001110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64110 - 64114

  --1111101001110011    1111101001110100    1111101001110101    1111101001110110    1111101001110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64115 - 64119

  --1111101001111000    1111101001111001    1111101001111010    1111101001111011    1111101001111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64120 - 64124

  --1111101001111101    1111101001111110    1111101001111111    1111101010000000    1111101010000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64125 - 64129

  --1111101010000010    1111101010000011    1111101010000100    1111101010000101    1111101010000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64130 - 64134

  --1111101010000111    1111101010001000    1111101010001001    1111101010001010    1111101010001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64135 - 64139

  --1111101010001100    1111101010001101    1111101010001110    1111101010001111    1111101010010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64140 - 64144

  --1111101010010001    1111101010010010    1111101010010011    1111101010010100    1111101010010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64145 - 64149

  --1111101010010110    1111101010010111    1111101010011000    1111101010011001    1111101010011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64150 - 64154

  --1111101010011011    1111101010011100    1111101010011101    1111101010011110    1111101010011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64155 - 64159

  --1111101010100000    1111101010100001    1111101010100010    1111101010100011    1111101010100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64160 - 64164

  --1111101010100101    1111101010100110    1111101010100111    1111101010101000    1111101010101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64165 - 64169

  --1111101010101010    1111101010101011    1111101010101100    1111101010101101    1111101010101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64170 - 64174

  --1111101010101111    1111101010110000    1111101010110001    1111101010110010    1111101010110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64175 - 64179

  --1111101010110100    1111101010110101    1111101010110110    1111101010110111    1111101010111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64180 - 64184

  --1111101010111001    1111101010111010    1111101010111011    1111101010111100    1111101010111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64185 - 64189

  --1111101010111110    1111101010111111    1111101011000000    1111101011000001    1111101011000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64190 - 64194

  --1111101011000011    1111101011000100    1111101011000101    1111101011000110    1111101011000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64195 - 64199

  --1111101011001000    1111101011001001    1111101011001010    1111101011001011    1111101011001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64200 - 64204

  --1111101011001101    1111101011001110    1111101011001111    1111101011010000    1111101011010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64205 - 64209

  --1111101011010010    1111101011010011    1111101011010100    1111101011010101    1111101011010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64210 - 64214

  --1111101011010111    1111101011011000    1111101011011001    1111101011011010    1111101011011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64215 - 64219

  --1111101011011100    1111101011011101    1111101011011110    1111101011011111    1111101011100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64220 - 64224

  --1111101011100001    1111101011100010    1111101011100011    1111101011100100    1111101011100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64225 - 64229

  --1111101011100110    1111101011100111    1111101011101000    1111101011101001    1111101011101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64230 - 64234

  --1111101011101011    1111101011101100    1111101011101101    1111101011101110    1111101011101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64235 - 64239

  --1111101011110000    1111101011110001    1111101011110010    1111101011110011    1111101011110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64240 - 64244

  --1111101011110101    1111101011110110    1111101011110111    1111101011111000    1111101011111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64245 - 64249

  --1111101011111010    1111101011111011    1111101011111100    1111101011111101    1111101011111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64250 - 64254

  --1111101011111111    1111101100000000    1111101100000001    1111101100000010    1111101100000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64255 - 64259

  --1111101100000100    1111101100000101    1111101100000110    1111101100000111    1111101100001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64260 - 64264

  --1111101100001001    1111101100001010    1111101100001011    1111101100001100    1111101100001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64265 - 64269

  --1111101100001110    1111101100001111    1111101100010000    1111101100010001    1111101100010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64270 - 64274

  --1111101100010011    1111101100010100    1111101100010101    1111101100010110    1111101100010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64275 - 64279

  --1111101100011000    1111101100011001    1111101100011010    1111101100011011    1111101100011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64280 - 64284

  --1111101100011101    1111101100011110    1111101100011111    1111101100100000    1111101100100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64285 - 64289

  --1111101100100010    1111101100100011    1111101100100100    1111101100100101    1111101100100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64290 - 64294

  --1111101100100111    1111101100101000    1111101100101001    1111101100101010    1111101100101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64295 - 64299

  --1111101100101100    1111101100101101    1111101100101110    1111101100101111    1111101100110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64300 - 64304

  --1111101100110001    1111101100110010    1111101100110011    1111101100110100    1111101100110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64305 - 64309

  --1111101100110110    1111101100110111    1111101100111000    1111101100111001    1111101100111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64310 - 64314

  --1111101100111011    1111101100111100    1111101100111101    1111101100111110    1111101100111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64315 - 64319

  --1111101101000000    1111101101000001    1111101101000010    1111101101000011    1111101101000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64320 - 64324

  --1111101101000101    1111101101000110    1111101101000111    1111101101001000    1111101101001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64325 - 64329

  --1111101101001010    1111101101001011    1111101101001100    1111101101001101    1111101101001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64330 - 64334

  --1111101101001111    1111101101010000    1111101101010001    1111101101010010    1111101101010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64335 - 64339

  --1111101101010100    1111101101010101    1111101101010110    1111101101010111    1111101101011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64340 - 64344

  --1111101101011001    1111101101011010    1111101101011011    1111101101011100    1111101101011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64345 - 64349

  --1111101101011110    1111101101011111    1111101101100000    1111101101100001    1111101101100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64350 - 64354

  --1111101101100011    1111101101100100    1111101101100101    1111101101100110    1111101101100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64355 - 64359

  --1111101101101000    1111101101101001    1111101101101010    1111101101101011    1111101101101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64360 - 64364

  --1111101101101101    1111101101101110    1111101101101111    1111101101110000    1111101101110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64365 - 64369

  --1111101101110010    1111101101110011    1111101101110100    1111101101110101    1111101101110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64370 - 64374

  --1111101101110111    1111101101111000    1111101101111001    1111101101111010    1111101101111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64375 - 64379

  --1111101101111100    1111101101111101    1111101101111110    1111101101111111    1111101110000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64380 - 64384

  --1111101110000001    1111101110000010    1111101110000011    1111101110000100    1111101110000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64385 - 64389

  --1111101110000110    1111101110000111    1111101110001000    1111101110001001    1111101110001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64390 - 64394

  --1111101110001011    1111101110001100    1111101110001101    1111101110001110    1111101110001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64395 - 64399

  --1111101110010000    1111101110010001    1111101110010010    1111101110010011    1111101110010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64400 - 64404

  --1111101110010101    1111101110010110    1111101110010111    1111101110011000    1111101110011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64405 - 64409

  --1111101110011010    1111101110011011    1111101110011100    1111101110011101    1111101110011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64410 - 64414

  --1111101110011111    1111101110100000    1111101110100001    1111101110100010    1111101110100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64415 - 64419

  --1111101110100100    1111101110100101    1111101110100110    1111101110100111    1111101110101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64420 - 64424

  --1111101110101001    1111101110101010    1111101110101011    1111101110101100    1111101110101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64425 - 64429

  --1111101110101110    1111101110101111    1111101110110000    1111101110110001    1111101110110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64430 - 64434

  --1111101110110011    1111101110110100    1111101110110101    1111101110110110    1111101110110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64435 - 64439

  --1111101110111000    1111101110111001    1111101110111010    1111101110111011    1111101110111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64440 - 64444

  --1111101110111101    1111101110111110    1111101110111111    1111101111000000    1111101111000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64445 - 64449

  --1111101111000010    1111101111000011    1111101111000100    1111101111000101    1111101111000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64450 - 64454

  --1111101111000111    1111101111001000    1111101111001001    1111101111001010    1111101111001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64455 - 64459

  --1111101111001100    1111101111001101    1111101111001110    1111101111001111    1111101111010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64460 - 64464

  --1111101111010001    1111101111010010    1111101111010011    1111101111010100    1111101111010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64465 - 64469

  --1111101111010110    1111101111010111    1111101111011000    1111101111011001    1111101111011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64470 - 64474

  --1111101111011011    1111101111011100    1111101111011101    1111101111011110    1111101111011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64475 - 64479

  --1111101111100000    1111101111100001    1111101111100010    1111101111100011    1111101111100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64480 - 64484

  --1111101111100101    1111101111100110    1111101111100111    1111101111101000    1111101111101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64485 - 64489

  --1111101111101010    1111101111101011    1111101111101100    1111101111101101    1111101111101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64490 - 64494

  --1111101111101111    1111101111110000    1111101111110001    1111101111110010    1111101111110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64495 - 64499

  --1111101111110100    1111101111110101    1111101111110110    1111101111110111    1111101111111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64500 - 64504

  --1111101111111001    1111101111111010    1111101111111011    1111101111111100    1111101111111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64505 - 64509

  --1111101111111110    1111101111111111    1111110000000000    1111110000000001    1111110000000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64510 - 64514

  --1111110000000011    1111110000000100    1111110000000101    1111110000000110    1111110000000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64515 - 64519

  --1111110000001000    1111110000001001    1111110000001010    1111110000001011    1111110000001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64520 - 64524

  --1111110000001101    1111110000001110    1111110000001111    1111110000010000    1111110000010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64525 - 64529

  --1111110000010010    1111110000010011    1111110000010100    1111110000010101    1111110000010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64530 - 64534

  --1111110000010111    1111110000011000    1111110000011001    1111110000011010    1111110000011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64535 - 64539

  --1111110000011100    1111110000011101    1111110000011110    1111110000011111    1111110000100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64540 - 64544

  --1111110000100001    1111110000100010    1111110000100011    1111110000100100    1111110000100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64545 - 64549

  --1111110000100110    1111110000100111    1111110000101000    1111110000101001    1111110000101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64550 - 64554

  --1111110000101011    1111110000101100    1111110000101101    1111110000101110    1111110000101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64555 - 64559

  --1111110000110000    1111110000110001    1111110000110010    1111110000110011    1111110000110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64560 - 64564

  --1111110000110101    1111110000110110    1111110000110111    1111110000111000    1111110000111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64565 - 64569

  --1111110000111010    1111110000111011    1111110000111100    1111110000111101    1111110000111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64570 - 64574

  --1111110000111111    1111110001000000    1111110001000001    1111110001000010    1111110001000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64575 - 64579

  --1111110001000100    1111110001000101    1111110001000110    1111110001000111    1111110001001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64580 - 64584

  --1111110001001001    1111110001001010    1111110001001011    1111110001001100    1111110001001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64585 - 64589

  --1111110001001110    1111110001001111    1111110001010000    1111110001010001    1111110001010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64590 - 64594

  --1111110001010011    1111110001010100    1111110001010101    1111110001010110    1111110001010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64595 - 64599

  --1111110001011000    1111110001011001    1111110001011010    1111110001011011    1111110001011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64600 - 64604

  --1111110001011101    1111110001011110    1111110001011111    1111110001100000    1111110001100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64605 - 64609

  --1111110001100010    1111110001100011    1111110001100100    1111110001100101    1111110001100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64610 - 64614

  --1111110001100111    1111110001101000    1111110001101001    1111110001101010    1111110001101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64615 - 64619

  --1111110001101100    1111110001101101    1111110001101110    1111110001101111    1111110001110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64620 - 64624

  --1111110001110001    1111110001110010    1111110001110011    1111110001110100    1111110001110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64625 - 64629

  --1111110001110110    1111110001110111    1111110001111000    1111110001111001    1111110001111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64630 - 64634

  --1111110001111011    1111110001111100    1111110001111101    1111110001111110    1111110001111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64635 - 64639

  --1111110010000000    1111110010000001    1111110010000010    1111110010000011    1111110010000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64640 - 64644

  --1111110010000101    1111110010000110    1111110010000111    1111110010001000    1111110010001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64645 - 64649

  --1111110010001010    1111110010001011    1111110010001100    1111110010001101    1111110010001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64650 - 64654

  --1111110010001111    1111110010010000    1111110010010001    1111110010010010    1111110010010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64655 - 64659

  --1111110010010100    1111110010010101    1111110010010110    1111110010010111    1111110010011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64660 - 64664

  --1111110010011001    1111110010011010    1111110010011011    1111110010011100    1111110010011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64665 - 64669

  --1111110010011110    1111110010011111    1111110010100000    1111110010100001    1111110010100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64670 - 64674

  --1111110010100011    1111110010100100    1111110010100101    1111110010100110    1111110010100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64675 - 64679

  --1111110010101000    1111110010101001    1111110010101010    1111110010101011    1111110010101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64680 - 64684

  --1111110010101101    1111110010101110    1111110010101111    1111110010110000    1111110010110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64685 - 64689

  --1111110010110010    1111110010110011    1111110010110100    1111110010110101    1111110010110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64690 - 64694

  --1111110010110111    1111110010111000    1111110010111001    1111110010111010    1111110010111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64695 - 64699

  --1111110010111100    1111110010111101    1111110010111110    1111110010111111    1111110011000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64700 - 64704

  --1111110011000001    1111110011000010    1111110011000011    1111110011000100    1111110011000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64705 - 64709

  --1111110011000110    1111110011000111    1111110011001000    1111110011001001    1111110011001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64710 - 64714

  --1111110011001011    1111110011001100    1111110011001101    1111110011001110    1111110011001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64715 - 64719

  --1111110011010000    1111110011010001    1111110011010010    1111110011010011    1111110011010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64720 - 64724

  --1111110011010101    1111110011010110    1111110011010111    1111110011011000    1111110011011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64725 - 64729

  --1111110011011010    1111110011011011    1111110011011100    1111110011011101    1111110011011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64730 - 64734

  --1111110011011111    1111110011100000    1111110011100001    1111110011100010    1111110011100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64735 - 64739

  --1111110011100100    1111110011100101    1111110011100110    1111110011100111    1111110011101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64740 - 64744

  --1111110011101001    1111110011101010    1111110011101011    1111110011101100    1111110011101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64745 - 64749

  --1111110011101110    1111110011101111    1111110011110000    1111110011110001    1111110011110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64750 - 64754

  --1111110011110011    1111110011110100    1111110011110101    1111110011110110    1111110011110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64755 - 64759

  --1111110011111000    1111110011111001    1111110011111010    1111110011111011    1111110011111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64760 - 64764

  --1111110011111101    1111110011111110    1111110011111111    1111110100000000    1111110100000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64765 - 64769

  --1111110100000010    1111110100000011    1111110100000100    1111110100000101    1111110100000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64770 - 64774

  --1111110100000111    1111110100001000    1111110100001001    1111110100001010    1111110100001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64775 - 64779

  --1111110100001100    1111110100001101    1111110100001110    1111110100001111    1111110100010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64780 - 64784

  --1111110100010001    1111110100010010    1111110100010011    1111110100010100    1111110100010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64785 - 64789

  --1111110100010110    1111110100010111    1111110100011000    1111110100011001    1111110100011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64790 - 64794

  --1111110100011011    1111110100011100    1111110100011101    1111110100011110    1111110100011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64795 - 64799

  --1111110100100000    1111110100100001    1111110100100010    1111110100100011    1111110100100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64800 - 64804

  --1111110100100101    1111110100100110    1111110100100111    1111110100101000    1111110100101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64805 - 64809

  --1111110100101010    1111110100101011    1111110100101100    1111110100101101    1111110100101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64810 - 64814

  --1111110100101111    1111110100110000    1111110100110001    1111110100110010    1111110100110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64815 - 64819

  --1111110100110100    1111110100110101    1111110100110110    1111110100110111    1111110100111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64820 - 64824

  --1111110100111001    1111110100111010    1111110100111011    1111110100111100    1111110100111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64825 - 64829

  --1111110100111110    1111110100111111    1111110101000000    1111110101000001    1111110101000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64830 - 64834

  --1111110101000011    1111110101000100    1111110101000101    1111110101000110    1111110101000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64835 - 64839

  --1111110101001000    1111110101001001    1111110101001010    1111110101001011    1111110101001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64840 - 64844

  --1111110101001101    1111110101001110    1111110101001111    1111110101010000    1111110101010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64845 - 64849

  --1111110101010010    1111110101010011    1111110101010100    1111110101010101    1111110101010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64850 - 64854

  --1111110101010111    1111110101011000    1111110101011001    1111110101011010    1111110101011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64855 - 64859

  --1111110101011100    1111110101011101    1111110101011110    1111110101011111    1111110101100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64860 - 64864

  --1111110101100001    1111110101100010    1111110101100011    1111110101100100    1111110101100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64865 - 64869

  --1111110101100110    1111110101100111    1111110101101000    1111110101101001    1111110101101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64870 - 64874

  --1111110101101011    1111110101101100    1111110101101101    1111110101101110    1111110101101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64875 - 64879

  --1111110101110000    1111110101110001    1111110101110010    1111110101110011    1111110101110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64880 - 64884

  --1111110101110101    1111110101110110    1111110101110111    1111110101111000    1111110101111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64885 - 64889

  --1111110101111010    1111110101111011    1111110101111100    1111110101111101    1111110101111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64890 - 64894

  --1111110101111111    1111110110000000    1111110110000001    1111110110000010    1111110110000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64895 - 64899

  --1111110110000100    1111110110000101    1111110110000110    1111110110000111    1111110110001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64900 - 64904

  --1111110110001001    1111110110001010    1111110110001011    1111110110001100    1111110110001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64905 - 64909

  --1111110110001110    1111110110001111    1111110110010000    1111110110010001    1111110110010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64910 - 64914

  --1111110110010011    1111110110010100    1111110110010101    1111110110010110    1111110110010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64915 - 64919

  --1111110110011000    1111110110011001    1111110110011010    1111110110011011    1111110110011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64920 - 64924

  --1111110110011101    1111110110011110    1111110110011111    1111110110100000    1111110110100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64925 - 64929

  --1111110110100010    1111110110100011    1111110110100100    1111110110100101    1111110110100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64930 - 64934

  --1111110110100111    1111110110101000    1111110110101001    1111110110101010    1111110110101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64935 - 64939

  --1111110110101100    1111110110101101    1111110110101110    1111110110101111    1111110110110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64940 - 64944

  --1111110110110001    1111110110110010    1111110110110011    1111110110110100    1111110110110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64945 - 64949

  --1111110110110110    1111110110110111    1111110110111000    1111110110111001    1111110110111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64950 - 64954

  --1111110110111011    1111110110111100    1111110110111101    1111110110111110    1111110110111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64955 - 64959

  --1111110111000000    1111110111000001    1111110111000010    1111110111000011    1111110111000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64960 - 64964

  --1111110111000101    1111110111000110    1111110111000111    1111110111001000    1111110111001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64965 - 64969

  --1111110111001010    1111110111001011    1111110111001100    1111110111001101    1111110111001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64970 - 64974

  --1111110111001111    1111110111010000    1111110111010001    1111110111010010    1111110111010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64975 - 64979

  --1111110111010100    1111110111010101    1111110111010110    1111110111010111    1111110111011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64980 - 64984

  --1111110111011001    1111110111011010    1111110111011011    1111110111011100    1111110111011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64985 - 64989

  --1111110111011110    1111110111011111    1111110111100000    1111110111100001    1111110111100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64990 - 64994

  --1111110111100011    1111110111100100    1111110111100101    1111110111100110    1111110111100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 64995 - 64999

  --1111110111101000    1111110111101001    1111110111101010    1111110111101011    1111110111101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65000 - 65004

  --1111110111101101    1111110111101110    1111110111101111    1111110111110000    1111110111110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65005 - 65009

  --1111110111110010    1111110111110011    1111110111110100    1111110111110101    1111110111110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65010 - 65014

  --1111110111110111    1111110111111000    1111110111111001    1111110111111010    1111110111111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65015 - 65019

  --1111110111111100    1111110111111101    1111110111111110    1111110111111111    1111111000000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65020 - 65024

  --1111111000000001    1111111000000010    1111111000000011    1111111000000100    1111111000000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65025 - 65029

  --1111111000000110    1111111000000111    1111111000001000    1111111000001001    1111111000001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65030 - 65034

  --1111111000001011    1111111000001100    1111111000001101    1111111000001110    1111111000001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65035 - 65039

  --1111111000010000    1111111000010001    1111111000010010    1111111000010011    1111111000010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65040 - 65044

  --1111111000010101    1111111000010110    1111111000010111    1111111000011000    1111111000011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65045 - 65049

  --1111111000011010    1111111000011011    1111111000011100    1111111000011101    1111111000011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65050 - 65054

  --1111111000011111    1111111000100000    1111111000100001    1111111000100010    1111111000100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65055 - 65059

  --1111111000100100    1111111000100101    1111111000100110    1111111000100111    1111111000101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65060 - 65064

  --1111111000101001    1111111000101010    1111111000101011    1111111000101100    1111111000101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65065 - 65069

  --1111111000101110    1111111000101111    1111111000110000    1111111000110001    1111111000110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65070 - 65074

  --1111111000110011    1111111000110100    1111111000110101    1111111000110110    1111111000110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65075 - 65079

  --1111111000111000    1111111000111001    1111111000111010    1111111000111011    1111111000111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65080 - 65084

  --1111111000111101    1111111000111110    1111111000111111    1111111001000000    1111111001000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65085 - 65089

  --1111111001000010    1111111001000011    1111111001000100    1111111001000101    1111111001000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65090 - 65094

  --1111111001000111    1111111001001000    1111111001001001    1111111001001010    1111111001001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65095 - 65099

  --1111111001001100    1111111001001101    1111111001001110    1111111001001111    1111111001010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65100 - 65104

  --1111111001010001    1111111001010010    1111111001010011    1111111001010100    1111111001010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65105 - 65109

  --1111111001010110    1111111001010111    1111111001011000    1111111001011001    1111111001011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65110 - 65114

  --1111111001011011    1111111001011100    1111111001011101    1111111001011110    1111111001011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65115 - 65119

  --1111111001100000    1111111001100001    1111111001100010    1111111001100011    1111111001100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65120 - 65124

  --1111111001100101    1111111001100110    1111111001100111    1111111001101000    1111111001101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65125 - 65129

  --1111111001101010    1111111001101011    1111111001101100    1111111001101101    1111111001101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65130 - 65134

  --1111111001101111    1111111001110000    1111111001110001    1111111001110010    1111111001110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65135 - 65139

  --1111111001110100    1111111001110101    1111111001110110    1111111001110111    1111111001111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65140 - 65144

  --1111111001111001    1111111001111010    1111111001111011    1111111001111100    1111111001111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65145 - 65149

  --1111111001111110    1111111001111111    1111111010000000    1111111010000001    1111111010000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65150 - 65154

  --1111111010000011    1111111010000100    1111111010000101    1111111010000110    1111111010000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65155 - 65159

  --1111111010001000    1111111010001001    1111111010001010    1111111010001011    1111111010001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65160 - 65164

  --1111111010001101    1111111010001110    1111111010001111    1111111010010000    1111111010010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65165 - 65169

  --1111111010010010    1111111010010011    1111111010010100    1111111010010101    1111111010010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65170 - 65174

  --1111111010010111    1111111010011000    1111111010011001    1111111010011010    1111111010011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65175 - 65179

  --1111111010011100    1111111010011101    1111111010011110    1111111010011111    1111111010100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65180 - 65184

  --1111111010100001    1111111010100010    1111111010100011    1111111010100100    1111111010100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65185 - 65189

  --1111111010100110    1111111010100111    1111111010101000    1111111010101001    1111111010101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65190 - 65194

  --1111111010101011    1111111010101100    1111111010101101    1111111010101110    1111111010101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65195 - 65199

  --1111111010110000    1111111010110001    1111111010110010    1111111010110011    1111111010110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65200 - 65204

  --1111111010110101    1111111010110110    1111111010110111    1111111010111000    1111111010111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65205 - 65209

  --1111111010111010    1111111010111011    1111111010111100    1111111010111101    1111111010111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65210 - 65214

  --1111111010111111    1111111011000000    1111111011000001    1111111011000010    1111111011000011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65215 - 65219

  --1111111011000100    1111111011000101    1111111011000110    1111111011000111    1111111011001000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65220 - 65224

  --1111111011001001    1111111011001010    1111111011001011    1111111011001100    1111111011001101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65225 - 65229

  --1111111011001110    1111111011001111    1111111011010000    1111111011010001    1111111011010010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65230 - 65234

  --1111111011010011    1111111011010100    1111111011010101    1111111011010110    1111111011010111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65235 - 65239

  --1111111011011000    1111111011011001    1111111011011010    1111111011011011    1111111011011100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65240 - 65244

  --1111111011011101    1111111011011110    1111111011011111    1111111011100000    1111111011100001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65245 - 65249

  --1111111011100010    1111111011100011    1111111011100100    1111111011100101    1111111011100110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65250 - 65254

  --1111111011100111    1111111011101000    1111111011101001    1111111011101010    1111111011101011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65255 - 65259

  --1111111011101100    1111111011101101    1111111011101110    1111111011101111    1111111011110000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65260 - 65264

  --1111111011110001    1111111011110010    1111111011110011    1111111011110100    1111111011110101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65265 - 65269

  --1111111011110110    1111111011110111    1111111011111000    1111111011111001    1111111011111010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65270 - 65274

  --1111111011111011    1111111011111100    1111111011111101    1111111011111110    1111111011111111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65275 - 65279

  --1111111100000000    1111111100000001    1111111100000010    1111111100000011    1111111100000100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65280 - 65284

  --1111111100000101    1111111100000110    1111111100000111    1111111100001000    1111111100001001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65285 - 65289

  --1111111100001010    1111111100001011    1111111100001100    1111111100001101    1111111100001110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65290 - 65294

  --1111111100001111    1111111100010000    1111111100010001    1111111100010010    1111111100010011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65295 - 65299

  --1111111100010100    1111111100010101    1111111100010110    1111111100010111    1111111100011000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65300 - 65304

  --1111111100011001    1111111100011010    1111111100011011    1111111100011100    1111111100011101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65305 - 65309

  --1111111100011110    1111111100011111    1111111100100000    1111111100100001    1111111100100010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65310 - 65314

  --1111111100100011    1111111100100100    1111111100100101    1111111100100110    1111111100100111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65315 - 65319

  --1111111100101000    1111111100101001    1111111100101010    1111111100101011    1111111100101100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65320 - 65324

  --1111111100101101    1111111100101110    1111111100101111    1111111100110000    1111111100110001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65325 - 65329

  --1111111100110010    1111111100110011    1111111100110100    1111111100110101    1111111100110110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65330 - 65334

  --1111111100110111    1111111100111000    1111111100111001    1111111100111010    1111111100111011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65335 - 65339

  --1111111100111100    1111111100111101    1111111100111110    1111111100111111    1111111101000000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65340 - 65344

  --1111111101000001    1111111101000010    1111111101000011    1111111101000100    1111111101000101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65345 - 65349

  --1111111101000110    1111111101000111    1111111101001000    1111111101001001    1111111101001010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65350 - 65354

  --1111111101001011    1111111101001100    1111111101001101    1111111101001110    1111111101001111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65355 - 65359

  --1111111101010000    1111111101010001    1111111101010010    1111111101010011    1111111101010100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65360 - 65364

  --1111111101010101    1111111101010110    1111111101010111    1111111101011000    1111111101011001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65365 - 65369

  --1111111101011010    1111111101011011    1111111101011100    1111111101011101    1111111101011110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65370 - 65374

  --1111111101011111    1111111101100000    1111111101100001    1111111101100010    1111111101100011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65375 - 65379

  --1111111101100100    1111111101100101    1111111101100110    1111111101100111    1111111101101000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65380 - 65384

  --1111111101101001    1111111101101010    1111111101101011    1111111101101100    1111111101101101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65385 - 65389

  --1111111101101110    1111111101101111    1111111101110000    1111111101110001    1111111101110010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65390 - 65394

  --1111111101110011    1111111101110100    1111111101110101    1111111101110110    1111111101110111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65395 - 65399

  --1111111101111000    1111111101111001    1111111101111010    1111111101111011    1111111101111100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65400 - 65404

  --1111111101111101    1111111101111110    1111111101111111    1111111110000000    1111111110000001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65405 - 65409

  --1111111110000010    1111111110000011    1111111110000100    1111111110000101    1111111110000110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65410 - 65414

  --1111111110000111    1111111110001000    1111111110001001    1111111110001010    1111111110001011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65415 - 65419

  --1111111110001100    1111111110001101    1111111110001110    1111111110001111    1111111110010000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65420 - 65424

  --1111111110010001    1111111110010010    1111111110010011    1111111110010100    1111111110010101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65425 - 65429

  --1111111110010110    1111111110010111    1111111110011000    1111111110011001    1111111110011010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65430 - 65434

  --1111111110011011    1111111110011100    1111111110011101    1111111110011110    1111111110011111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65435 - 65439

  --1111111110100000    1111111110100001    1111111110100010    1111111110100011    1111111110100100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65440 - 65444

  --1111111110100101    1111111110100110    1111111110100111    1111111110101000    1111111110101001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65445 - 65449

  --1111111110101010    1111111110101011    1111111110101100    1111111110101101    1111111110101110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65450 - 65454

  --1111111110101111    1111111110110000    1111111110110001    1111111110110010    1111111110110011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65455 - 65459

  --1111111110110100    1111111110110101    1111111110110110    1111111110110111    1111111110111000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65460 - 65464

  --1111111110111001    1111111110111010    1111111110111011    1111111110111100    1111111110111101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65465 - 65469

  --1111111110111110    1111111110111111    1111111111000000    1111111111000001    1111111111000010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65470 - 65474

  --1111111111000011    1111111111000100    1111111111000101    1111111111000110    1111111111000111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65475 - 65479

  --1111111111001000    1111111111001001    1111111111001010    1111111111001011    1111111111001100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65480 - 65484

  --1111111111001101    1111111111001110    1111111111001111    1111111111010000    1111111111010001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65485 - 65489

  --1111111111010010    1111111111010011    1111111111010100    1111111111010101    1111111111010110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65490 - 65494

  --1111111111010111    1111111111011000    1111111111011001    1111111111011010    1111111111011011    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65495 - 65499

  --1111111111011100    1111111111011101    1111111111011110    1111111111011111    1111111111100000    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65500 - 65504

  --1111111111100001    1111111111100010    1111111111100011    1111111111100100    1111111111100101    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65505 - 65509

  --1111111111100110    1111111111100111    1111111111101000    1111111111101001    1111111111101010    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65510 - 65514

  --1111111111101011    1111111111101100    1111111111101101    1111111111101110    1111111111101111    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65515 - 65519

  --1111111111110000    1111111111110001    1111111111110010    1111111111110011    1111111111110100    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65520 - 65524

  --1111111111110101    1111111111110110    1111111111110111    1111111111111000    1111111111111001    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65525 - 65529

  --1111111111111010    1111111111111011    1111111111111100    1111111111111101    1111111111111110    
   "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", -- 65530 - 65534

  --1111111111111111 
   "0000000000000000"										       															 -- 65535

	);
	
begin
	
	data <= rom(to_integer(unsigned(address)));

end architecture;
	